
// 	Fri Dec 23 14:10:30 2022
//	vlsi
//	localhost.localdomain

module registerNbits (clk_CTS_0_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits

module registerNbits__0_9 (clk_CTS_0_PP_0, clk_CTS_0_PP_1, clk_CTS_0_PP_2, clk, reset, 
    en, inp, out);

output [31:0] out;
output clk_CTS_0_PP_0;
output clk_CTS_0_PP_1;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_2;
wire n_0_0;
wire n_1;
wire CTS_n_tid0_25;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid0_34;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X2 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid0_25), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid0_25), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid0_25), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid0_25), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid0_25), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid0_25), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid0_25), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid0_25), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid0_25), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid0_25), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid0_25), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid0_25), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid0_25), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid0_25), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid0_25), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid0_25), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid0_25), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid0_25), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid0_25), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid0_25), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid0_25), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid0_25), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid0_25), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid0_25), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid0_25), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid0_25), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid0_25), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid0_25), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid0_25), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid0_25), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid0_25), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid0_25), .D (n_33));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n_tid0_25), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
INV_X4 CTS_L3_c_tid0_29 (.ZN (clk_CTS_0_PP_1), .A (CTS_n_tid0_34));
CLKBUF_X3 CTS_L4_c_tid0_27 (.Z (clk_CTS_0_PP_0), .A (clk_CTS_0_PP_1));
INV_X8 CTS_L2_c_tid0_30 (.ZN (CTS_n_tid0_34), .A (clk_CTS_0_PP_2));

endmodule //registerNbits__0_9

module datapath (inputB, inputA, result);

output [63:0] result;
input [31:0] inputA;
input [31:0] inputB;
wire n_2985;
wire n_3397;
wire n_1;
wire n_0;
wire n_2955;
wire n_2984;
wire n_3013;
wire n_3;
wire n_2;
wire n_3041;
wire n_5;
wire n_4;
wire n_2925;
wire n_2954;
wire n_2983;
wire n_7;
wire n_6;
wire n_3012;
wire n_3040;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_2896;
wire n_2924;
wire n_2953;
wire n_13;
wire n_12;
wire n_2982;
wire n_3011;
wire n_3039;
wire n_15;
wire n_14;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_2865;
wire n_2895;
wire n_2923;
wire n_21;
wire n_20;
wire n_2952;
wire n_2981;
wire n_3010;
wire n_23;
wire n_22;
wire n_3038;
wire n_25;
wire n_24;
wire n_27;
wire n_26;
wire n_29;
wire n_28;
wire n_2835;
wire n_2864;
wire n_2894;
wire n_31;
wire n_30;
wire n_2922;
wire n_2951;
wire n_2980;
wire n_33;
wire n_32;
wire n_3009;
wire n_3037;
wire n_35;
wire n_34;
wire n_37;
wire n_36;
wire n_39;
wire n_38;
wire n_41;
wire n_40;
wire n_2806;
wire n_2834;
wire n_2863;
wire n_43;
wire n_42;
wire n_2893;
wire n_2921;
wire n_2950;
wire n_45;
wire n_44;
wire n_2979;
wire n_3008;
wire n_3036;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_53;
wire n_52;
wire n_55;
wire n_54;
wire n_2775;
wire n_2805;
wire n_2833;
wire n_57;
wire n_56;
wire n_2862;
wire n_2892;
wire n_2920;
wire n_59;
wire n_58;
wire n_2949;
wire n_2978;
wire n_3007;
wire n_61;
wire n_60;
wire n_3035;
wire n_63;
wire n_62;
wire n_65;
wire n_64;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_71;
wire n_70;
wire n_2745;
wire n_2774;
wire n_2804;
wire n_73;
wire n_72;
wire n_2832;
wire n_2861;
wire n_2891;
wire n_75;
wire n_74;
wire n_2919;
wire n_2948;
wire n_2977;
wire n_77;
wire n_76;
wire n_3006;
wire n_3034;
wire n_79;
wire n_78;
wire n_81;
wire n_80;
wire n_83;
wire n_82;
wire n_85;
wire n_84;
wire n_87;
wire n_86;
wire n_89;
wire n_88;
wire n_2716;
wire n_2744;
wire n_2773;
wire n_91;
wire n_90;
wire n_2803;
wire n_2831;
wire n_2860;
wire n_93;
wire n_92;
wire n_2890;
wire n_2918;
wire n_2947;
wire n_95;
wire n_94;
wire n_2976;
wire n_3005;
wire n_3033;
wire n_97;
wire n_96;
wire n_99;
wire n_98;
wire n_101;
wire n_100;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_107;
wire n_106;
wire n_109;
wire n_108;
wire n_2685;
wire n_2715;
wire n_2743;
wire n_111;
wire n_110;
wire n_2772;
wire n_2802;
wire n_2830;
wire n_113;
wire n_112;
wire n_2859;
wire n_2889;
wire n_2917;
wire n_115;
wire n_114;
wire n_2946;
wire n_2975;
wire n_3004;
wire n_117;
wire n_116;
wire n_3032;
wire n_119;
wire n_118;
wire n_121;
wire n_120;
wire n_123;
wire n_122;
wire n_125;
wire n_124;
wire n_127;
wire n_126;
wire n_129;
wire n_128;
wire n_131;
wire n_130;
wire n_2655;
wire n_2684;
wire n_2714;
wire n_133;
wire n_132;
wire n_2742;
wire n_2771;
wire n_2801;
wire n_135;
wire n_134;
wire n_2829;
wire n_2858;
wire n_2888;
wire n_137;
wire n_136;
wire n_2916;
wire n_2945;
wire n_2974;
wire n_139;
wire n_138;
wire n_3003;
wire n_3031;
wire n_141;
wire n_140;
wire n_143;
wire n_142;
wire n_145;
wire n_144;
wire n_147;
wire n_146;
wire n_149;
wire n_148;
wire n_151;
wire n_150;
wire n_153;
wire n_152;
wire n_155;
wire n_154;
wire n_2626;
wire n_2654;
wire n_2683;
wire n_157;
wire n_156;
wire n_2713;
wire n_2741;
wire n_2770;
wire n_159;
wire n_158;
wire n_2800;
wire n_2828;
wire n_2857;
wire n_161;
wire n_160;
wire n_2887;
wire n_2915;
wire n_2944;
wire n_163;
wire n_162;
wire n_2973;
wire n_3002;
wire n_3030;
wire n_165;
wire n_164;
wire n_167;
wire n_166;
wire n_169;
wire n_168;
wire n_171;
wire n_170;
wire n_173;
wire n_172;
wire n_175;
wire n_174;
wire n_177;
wire n_176;
wire n_179;
wire n_178;
wire n_181;
wire n_180;
wire n_2595;
wire n_2625;
wire n_2653;
wire n_183;
wire n_182;
wire n_2682;
wire n_2712;
wire n_2740;
wire n_185;
wire n_184;
wire n_2769;
wire n_2799;
wire n_2827;
wire n_187;
wire n_186;
wire n_2856;
wire n_2886;
wire n_2914;
wire n_189;
wire n_188;
wire n_2943;
wire n_2972;
wire n_3001;
wire n_191;
wire n_190;
wire n_3029;
wire n_193;
wire n_192;
wire n_195;
wire n_194;
wire n_197;
wire n_196;
wire n_199;
wire n_198;
wire n_201;
wire n_200;
wire n_203;
wire n_202;
wire n_205;
wire n_204;
wire n_207;
wire n_206;
wire n_209;
wire n_208;
wire n_2565;
wire n_2594;
wire n_2624;
wire n_211;
wire n_210;
wire n_2652;
wire n_2681;
wire n_2711;
wire n_213;
wire n_212;
wire n_2739;
wire n_2768;
wire n_2798;
wire n_215;
wire n_214;
wire n_2826;
wire n_2855;
wire n_2885;
wire n_217;
wire n_216;
wire n_2913;
wire n_2942;
wire n_2971;
wire n_219;
wire n_218;
wire n_3000;
wire n_3028;
wire n_221;
wire n_220;
wire n_223;
wire n_222;
wire n_225;
wire n_224;
wire n_227;
wire n_226;
wire n_229;
wire n_228;
wire n_231;
wire n_230;
wire n_233;
wire n_232;
wire n_235;
wire n_234;
wire n_237;
wire n_236;
wire n_239;
wire n_238;
wire n_2536;
wire n_2564;
wire n_2593;
wire n_241;
wire n_240;
wire n_2623;
wire n_2651;
wire n_2680;
wire n_243;
wire n_242;
wire n_2710;
wire n_2738;
wire n_2767;
wire n_245;
wire n_244;
wire n_2797;
wire n_2825;
wire n_2854;
wire n_247;
wire n_246;
wire n_2884;
wire n_2912;
wire n_2941;
wire n_249;
wire n_248;
wire n_2970;
wire n_2999;
wire n_3027;
wire n_251;
wire n_250;
wire n_253;
wire n_252;
wire n_255;
wire n_254;
wire n_257;
wire n_256;
wire n_259;
wire n_258;
wire n_261;
wire n_260;
wire n_263;
wire n_262;
wire n_265;
wire n_264;
wire n_267;
wire n_266;
wire n_269;
wire n_268;
wire n_271;
wire n_270;
wire n_2505;
wire n_2535;
wire n_2563;
wire n_273;
wire n_272;
wire n_2592;
wire n_2622;
wire n_2650;
wire n_275;
wire n_274;
wire n_2679;
wire n_2709;
wire n_2737;
wire n_277;
wire n_276;
wire n_2766;
wire n_2796;
wire n_2824;
wire n_279;
wire n_278;
wire n_2853;
wire n_2883;
wire n_2911;
wire n_281;
wire n_280;
wire n_2940;
wire n_2969;
wire n_2998;
wire n_283;
wire n_282;
wire n_3026;
wire n_285;
wire n_284;
wire n_287;
wire n_286;
wire n_289;
wire n_288;
wire n_291;
wire n_290;
wire n_293;
wire n_292;
wire n_295;
wire n_294;
wire n_297;
wire n_296;
wire n_299;
wire n_298;
wire n_301;
wire n_300;
wire n_303;
wire n_302;
wire n_305;
wire n_304;
wire n_2475;
wire n_2504;
wire n_2534;
wire n_307;
wire n_306;
wire n_2562;
wire n_2591;
wire n_2621;
wire n_309;
wire n_308;
wire n_2649;
wire n_2678;
wire n_2708;
wire n_311;
wire n_310;
wire n_2736;
wire n_2765;
wire n_2795;
wire n_313;
wire n_312;
wire n_2823;
wire n_2852;
wire n_2882;
wire n_315;
wire n_314;
wire n_2910;
wire n_2939;
wire n_2968;
wire n_317;
wire n_316;
wire n_2997;
wire n_3025;
wire n_319;
wire n_318;
wire n_321;
wire n_320;
wire n_323;
wire n_322;
wire n_325;
wire n_324;
wire n_327;
wire n_326;
wire n_329;
wire n_328;
wire n_331;
wire n_330;
wire n_333;
wire n_332;
wire n_335;
wire n_334;
wire n_337;
wire n_336;
wire n_339;
wire n_338;
wire n_341;
wire n_340;
wire n_2446;
wire n_2474;
wire n_2503;
wire n_343;
wire n_342;
wire n_2533;
wire n_2561;
wire n_2590;
wire n_345;
wire n_344;
wire n_2620;
wire n_2648;
wire n_2677;
wire n_347;
wire n_346;
wire n_2707;
wire n_2735;
wire n_2764;
wire n_349;
wire n_348;
wire n_2794;
wire n_2822;
wire n_2851;
wire n_351;
wire n_350;
wire n_2881;
wire n_2909;
wire n_2938;
wire n_353;
wire n_352;
wire n_2967;
wire n_2996;
wire n_3024;
wire n_355;
wire n_354;
wire n_357;
wire n_356;
wire n_359;
wire n_358;
wire n_361;
wire n_360;
wire n_363;
wire n_362;
wire n_365;
wire n_364;
wire n_367;
wire n_366;
wire n_369;
wire n_368;
wire n_371;
wire n_370;
wire n_373;
wire n_372;
wire n_375;
wire n_374;
wire n_377;
wire n_376;
wire n_379;
wire n_378;
wire n_2415;
wire n_2445;
wire n_2473;
wire n_381;
wire n_380;
wire n_2502;
wire n_2532;
wire n_2560;
wire n_383;
wire n_382;
wire n_2589;
wire n_2619;
wire n_2647;
wire n_385;
wire n_384;
wire n_2676;
wire n_2706;
wire n_2734;
wire n_387;
wire n_386;
wire n_2763;
wire n_2793;
wire n_2821;
wire n_389;
wire n_388;
wire n_2850;
wire n_2880;
wire n_2908;
wire n_391;
wire n_390;
wire n_2937;
wire n_2966;
wire n_2995;
wire n_393;
wire n_392;
wire n_3023;
wire n_395;
wire n_394;
wire n_397;
wire n_396;
wire n_399;
wire n_398;
wire n_401;
wire n_400;
wire n_403;
wire n_402;
wire n_405;
wire n_404;
wire n_407;
wire n_406;
wire n_409;
wire n_408;
wire n_411;
wire n_410;
wire n_413;
wire n_412;
wire n_415;
wire n_414;
wire n_417;
wire n_416;
wire n_419;
wire n_418;
wire n_2385;
wire n_2414;
wire n_2444;
wire n_421;
wire n_420;
wire n_2472;
wire n_2501;
wire n_2531;
wire n_423;
wire n_422;
wire n_2559;
wire n_2588;
wire n_2618;
wire n_425;
wire n_424;
wire n_2646;
wire n_2675;
wire n_2705;
wire n_427;
wire n_426;
wire n_2733;
wire n_2762;
wire n_2792;
wire n_429;
wire n_428;
wire n_2820;
wire n_2849;
wire n_2879;
wire n_431;
wire n_430;
wire n_2907;
wire n_2936;
wire n_2965;
wire n_433;
wire n_432;
wire n_2994;
wire n_3022;
wire n_435;
wire n_434;
wire n_437;
wire n_436;
wire n_439;
wire n_438;
wire n_441;
wire n_440;
wire n_443;
wire n_442;
wire n_445;
wire n_444;
wire n_447;
wire n_446;
wire n_449;
wire n_448;
wire n_451;
wire n_450;
wire n_453;
wire n_452;
wire n_455;
wire n_454;
wire n_457;
wire n_456;
wire n_459;
wire n_458;
wire n_461;
wire n_460;
wire n_2356;
wire n_2384;
wire n_2413;
wire n_463;
wire n_462;
wire n_2443;
wire n_2471;
wire n_2500;
wire n_465;
wire n_464;
wire n_2530;
wire n_2558;
wire n_2587;
wire n_467;
wire n_466;
wire n_2617;
wire n_2645;
wire n_2674;
wire n_469;
wire n_468;
wire n_2704;
wire n_2732;
wire n_2761;
wire n_471;
wire n_470;
wire n_2791;
wire n_2819;
wire n_2848;
wire n_473;
wire n_472;
wire n_2878;
wire n_2906;
wire n_2935;
wire n_475;
wire n_474;
wire n_2964;
wire n_2993;
wire n_3021;
wire n_477;
wire n_476;
wire n_479;
wire n_478;
wire n_481;
wire n_480;
wire n_483;
wire n_482;
wire n_485;
wire n_484;
wire n_487;
wire n_486;
wire n_489;
wire n_488;
wire n_491;
wire n_490;
wire n_493;
wire n_492;
wire n_495;
wire n_494;
wire n_497;
wire n_496;
wire n_499;
wire n_498;
wire n_501;
wire n_500;
wire n_503;
wire n_502;
wire n_505;
wire n_504;
wire n_2325;
wire n_2355;
wire n_2383;
wire n_507;
wire n_506;
wire n_2412;
wire n_2442;
wire n_2470;
wire n_509;
wire n_508;
wire n_2499;
wire n_2529;
wire n_2557;
wire n_511;
wire n_510;
wire n_2586;
wire n_2616;
wire n_2644;
wire n_513;
wire n_512;
wire n_2673;
wire n_2703;
wire n_2731;
wire n_515;
wire n_514;
wire n_2760;
wire n_2790;
wire n_2818;
wire n_517;
wire n_516;
wire n_2847;
wire n_2877;
wire n_2905;
wire n_519;
wire n_518;
wire n_2934;
wire n_2963;
wire n_2992;
wire n_521;
wire n_520;
wire n_3020;
wire n_523;
wire n_522;
wire n_525;
wire n_524;
wire n_527;
wire n_526;
wire n_529;
wire n_528;
wire n_531;
wire n_530;
wire n_533;
wire n_532;
wire n_535;
wire n_534;
wire n_537;
wire n_536;
wire n_539;
wire n_538;
wire n_541;
wire n_540;
wire n_543;
wire n_542;
wire n_545;
wire n_544;
wire n_547;
wire n_546;
wire n_549;
wire n_548;
wire n_551;
wire n_550;
wire n_2295;
wire n_2324;
wire n_2354;
wire n_553;
wire n_552;
wire n_2382;
wire n_2411;
wire n_2441;
wire n_555;
wire n_554;
wire n_2469;
wire n_2498;
wire n_2528;
wire n_557;
wire n_556;
wire n_2556;
wire n_2585;
wire n_2615;
wire n_559;
wire n_558;
wire n_2643;
wire n_2672;
wire n_2702;
wire n_561;
wire n_560;
wire n_2730;
wire n_2759;
wire n_2789;
wire n_563;
wire n_562;
wire n_2817;
wire n_2846;
wire n_2876;
wire n_565;
wire n_564;
wire n_2904;
wire n_2933;
wire n_2962;
wire n_567;
wire n_566;
wire n_2991;
wire n_3019;
wire n_569;
wire n_568;
wire n_571;
wire n_570;
wire n_573;
wire n_572;
wire n_575;
wire n_574;
wire n_577;
wire n_576;
wire n_579;
wire n_578;
wire n_581;
wire n_580;
wire n_583;
wire n_582;
wire n_585;
wire n_584;
wire n_587;
wire n_586;
wire n_589;
wire n_588;
wire n_591;
wire n_590;
wire n_593;
wire n_592;
wire n_595;
wire n_594;
wire n_597;
wire n_596;
wire n_599;
wire n_598;
wire n_2266;
wire n_2294;
wire n_2323;
wire n_601;
wire n_600;
wire n_2353;
wire n_2381;
wire n_2410;
wire n_603;
wire n_602;
wire n_2440;
wire n_2468;
wire n_2497;
wire n_605;
wire n_604;
wire n_2527;
wire n_2555;
wire n_2584;
wire n_607;
wire n_606;
wire n_2614;
wire n_2642;
wire n_2671;
wire n_609;
wire n_608;
wire n_2701;
wire n_2729;
wire n_2758;
wire n_611;
wire n_610;
wire n_2788;
wire n_2816;
wire n_2845;
wire n_613;
wire n_612;
wire n_2875;
wire n_2903;
wire n_2932;
wire n_615;
wire n_614;
wire n_2961;
wire n_2990;
wire n_3018;
wire n_617;
wire n_616;
wire n_619;
wire n_618;
wire n_621;
wire n_620;
wire n_623;
wire n_622;
wire n_625;
wire n_624;
wire n_627;
wire n_626;
wire n_629;
wire n_628;
wire n_631;
wire n_630;
wire n_633;
wire n_632;
wire n_635;
wire n_634;
wire n_637;
wire n_636;
wire n_639;
wire n_638;
wire n_641;
wire n_640;
wire n_643;
wire n_642;
wire n_645;
wire n_644;
wire n_647;
wire n_646;
wire n_649;
wire n_648;
wire n_2235;
wire n_2265;
wire n_2293;
wire n_651;
wire n_650;
wire n_2322;
wire n_2352;
wire n_2380;
wire n_653;
wire n_652;
wire n_2409;
wire n_2439;
wire n_2467;
wire n_655;
wire n_654;
wire n_2496;
wire n_2526;
wire n_2554;
wire n_657;
wire n_656;
wire n_2583;
wire n_2613;
wire n_2641;
wire n_659;
wire n_658;
wire n_2670;
wire n_2700;
wire n_2728;
wire n_661;
wire n_660;
wire n_2757;
wire n_2787;
wire n_2815;
wire n_663;
wire n_662;
wire n_2844;
wire n_2874;
wire n_2902;
wire n_665;
wire n_664;
wire n_2931;
wire n_2960;
wire n_2989;
wire n_667;
wire n_666;
wire n_3017;
wire n_669;
wire n_668;
wire n_671;
wire n_670;
wire n_673;
wire n_672;
wire n_675;
wire n_674;
wire n_677;
wire n_676;
wire n_679;
wire n_678;
wire n_681;
wire n_680;
wire n_683;
wire n_682;
wire n_685;
wire n_684;
wire n_687;
wire n_686;
wire n_689;
wire n_688;
wire n_691;
wire n_690;
wire n_693;
wire n_692;
wire n_695;
wire n_694;
wire n_697;
wire n_696;
wire n_699;
wire n_698;
wire n_701;
wire n_700;
wire n_2205;
wire n_2234;
wire n_2264;
wire n_703;
wire n_702;
wire n_2292;
wire n_2321;
wire n_2351;
wire n_705;
wire n_704;
wire n_2379;
wire n_2408;
wire n_2438;
wire n_707;
wire n_706;
wire n_2466;
wire n_2495;
wire n_2525;
wire n_709;
wire n_708;
wire n_2553;
wire n_2582;
wire n_2612;
wire n_711;
wire n_710;
wire n_2640;
wire n_2669;
wire n_2699;
wire n_713;
wire n_712;
wire n_2727;
wire n_2756;
wire n_2786;
wire n_715;
wire n_714;
wire n_2814;
wire n_2843;
wire n_2873;
wire n_717;
wire n_716;
wire n_2901;
wire n_2930;
wire n_2959;
wire n_719;
wire n_718;
wire n_2988;
wire n_3016;
wire n_721;
wire n_720;
wire n_723;
wire n_722;
wire n_725;
wire n_724;
wire n_727;
wire n_726;
wire n_729;
wire n_728;
wire n_731;
wire n_730;
wire n_733;
wire n_732;
wire n_735;
wire n_734;
wire n_737;
wire n_736;
wire n_739;
wire n_738;
wire n_741;
wire n_740;
wire n_743;
wire n_742;
wire n_745;
wire n_744;
wire n_747;
wire n_746;
wire n_749;
wire n_748;
wire n_751;
wire n_750;
wire n_753;
wire n_752;
wire n_755;
wire n_754;
wire n_2176;
wire n_2204;
wire n_2233;
wire n_757;
wire n_756;
wire n_2263;
wire n_2291;
wire n_2320;
wire n_759;
wire n_758;
wire n_777;
wire n_776;
wire n_779;
wire n_778;
wire n_781;
wire n_780;
wire n_783;
wire n_782;
wire n_898;
wire n_900;
wire n_870;
wire n_785;
wire n_784;
wire n_884;
wire n_886;
wire n_831;
wire n_787;
wire n_786;
wire n_832;
wire n_834;
wire n_789;
wire n_788;
wire n_791;
wire n_790;
wire n_793;
wire n_792;
wire n_795;
wire n_794;
wire n_797;
wire n_796;
wire n_799;
wire n_798;
wire n_801;
wire n_800;
wire n_803;
wire n_802;
wire n_805;
wire n_804;
wire n_807;
wire n_806;
wire n_809;
wire n_808;
wire n_811;
wire n_810;
wire n_2173;
wire n_2175;
wire n_2203;
wire n_813;
wire n_812;
wire n_2232;
wire n_2262;
wire n_2290;
wire n_815;
wire n_814;
wire n_2319;
wire n_2349;
wire n_2377;
wire n_817;
wire n_816;
wire n_2406;
wire n_2436;
wire n_2464;
wire n_819;
wire n_818;
wire n_2493;
wire n_2523;
wire n_2551;
wire n_821;
wire n_820;
wire n_2580;
wire n_2610;
wire n_2638;
wire n_823;
wire n_822;
wire n_2667;
wire n_2697;
wire n_2725;
wire n_825;
wire n_824;
wire n_2754;
wire n_2784;
wire n_2812;
wire n_827;
wire n_826;
wire n_2841;
wire n_2871;
wire n_2899;
wire n_829;
wire n_828;
wire n_839;
wire n_838;
wire n_982;
wire n_841;
wire n_840;
wire n_843;
wire n_842;
wire n_845;
wire n_844;
wire n_847;
wire n_846;
wire n_836;
wire n_849;
wire n_848;
wire n_894;
wire n_937;
wire n_851;
wire n_850;
wire n_853;
wire n_852;
wire n_855;
wire n_854;
wire n_857;
wire n_856;
wire n_859;
wire n_858;
wire n_861;
wire n_860;
wire n_863;
wire n_862;
wire n_865;
wire n_864;
wire n_867;
wire n_866;
wire n_869;
wire n_868;
wire n_889;
wire n_888;
wire n_891;
wire n_890;
wire n_893;
wire n_892;
wire n_2159;
wire n_1007;
wire n_770;
wire n_897;
wire n_896;
wire n_760;
wire n_2167;
wire n_903;
wire n_902;
wire n_905;
wire n_904;
wire n_907;
wire n_906;
wire n_939;
wire n_909;
wire n_908;
wire n_772;
wire n_911;
wire n_910;
wire n_774;
wire n_913;
wire n_912;
wire n_915;
wire n_914;
wire n_917;
wire n_916;
wire n_919;
wire n_918;
wire n_921;
wire n_920;
wire n_923;
wire n_922;
wire n_925;
wire n_924;
wire n_2174;
wire n_2201;
wire n_2230;
wire n_927;
wire n_926;
wire n_2260;
wire n_2288;
wire n_2317;
wire n_929;
wire n_928;
wire n_2347;
wire n_2375;
wire n_2404;
wire n_931;
wire n_930;
wire n_2434;
wire n_2462;
wire n_2491;
wire n_933;
wire n_932;
wire n_2521;
wire n_2549;
wire n_2578;
wire n_935;
wire n_934;
wire n_951;
wire n_950;
wire n_957;
wire n_956;
wire n_2153;
wire n_959;
wire n_958;
wire n_965;
wire n_964;
wire n_967;
wire n_966;
wire n_962;
wire n_1020;
wire n_969;
wire n_968;
wire n_830;
wire n_941;
wire n_971;
wire n_970;
wire n_973;
wire n_972;
wire n_975;
wire n_974;
wire n_977;
wire n_976;
wire n_979;
wire n_978;
wire n_981;
wire n_980;
wire n_2374;
wire n_2403;
wire n_2433;
wire n_987;
wire n_986;
wire n_2461;
wire n_2490;
wire n_2520;
wire n_989;
wire n_988;
wire n_2548;
wire n_2577;
wire n_2607;
wire n_991;
wire n_990;
wire n_2635;
wire n_2664;
wire n_2694;
wire n_993;
wire n_992;
wire n_2722;
wire n_2751;
wire n_2781;
wire n_995;
wire n_994;
wire n_2809;
wire n_2838;
wire n_2868;
wire n_997;
wire n_996;
wire n_1018;
wire n_952;
wire n_954;
wire n_999;
wire n_998;
wire n_960;
wire n_1001;
wire n_1000;
wire n_1003;
wire n_1002;
wire n_1009;
wire n_1008;
wire n_1011;
wire n_1010;
wire n_762;
wire n_764;
wire n_2139;
wire n_1013;
wire n_1012;
wire n_1015;
wire n_1014;
wire n_1017;
wire n_1016;
wire n_1023;
wire n_1022;
wire n_1067;
wire n_1025;
wire n_1024;
wire n_1027;
wire n_1026;
wire n_943;
wire n_1029;
wire n_1028;
wire n_1031;
wire n_1030;
wire n_1033;
wire n_1032;
wire n_1035;
wire n_1034;
wire n_2199;
wire n_2228;
wire n_2258;
wire n_1037;
wire n_1036;
wire n_2286;
wire n_2315;
wire n_2345;
wire n_1039;
wire n_1038;
wire n_2373;
wire n_2402;
wire n_2432;
wire n_1041;
wire n_1040;
wire n_2460;
wire n_2489;
wire n_2519;
wire n_1043;
wire n_1042;
wire n_2547;
wire n_2576;
wire n_2606;
wire n_1045;
wire n_1044;
wire n_2634;
wire n_2663;
wire n_2693;
wire n_1047;
wire n_1046;
wire n_2721;
wire n_2750;
wire n_2780;
wire n_1049;
wire n_1048;
wire n_2808;
wire n_2837;
wire n_2867;
wire n_1051;
wire n_1050;
wire n_1053;
wire n_1052;
wire n_1055;
wire n_1054;
wire n_1059;
wire n_1058;
wire n_2116;
wire n_1061;
wire n_1060;
wire n_1063;
wire n_1062;
wire n_1065;
wire n_1064;
wire n_1069;
wire n_1068;
wire n_1057;
wire n_1071;
wire n_1070;
wire n_1073;
wire n_1072;
wire n_1075;
wire n_1074;
wire n_1079;
wire n_1078;
wire n_1081;
wire n_1080;
wire n_1076;
wire n_1083;
wire n_1082;
wire n_1085;
wire n_1084;
wire n_1087;
wire n_1086;
wire n_2198;
wire n_2227;
wire n_2257;
wire n_1089;
wire n_1088;
wire n_2285;
wire n_2314;
wire n_2344;
wire n_1091;
wire n_1090;
wire n_2372;
wire n_2401;
wire n_2431;
wire n_1093;
wire n_1092;
wire n_2459;
wire n_2488;
wire n_2518;
wire n_1095;
wire n_1094;
wire n_2546;
wire n_2575;
wire n_2605;
wire n_1097;
wire n_1096;
wire n_2633;
wire n_2662;
wire n_2692;
wire n_1099;
wire n_1098;
wire n_2720;
wire n_2749;
wire n_2779;
wire n_1101;
wire n_1100;
wire n_2807;
wire n_2836;
wire n_2866;
wire n_1103;
wire n_1102;
wire n_1105;
wire n_1104;
wire n_1107;
wire n_1106;
wire n_2122;
wire n_766;
wire n_1109;
wire n_1108;
wire n_2115;
wire n_1111;
wire n_1110;
wire n_1113;
wire n_1112;
wire n_1115;
wire n_1114;
wire n_2109;
wire n_1117;
wire n_1116;
wire n_2102;
wire n_1119;
wire n_1118;
wire n_1121;
wire n_1120;
wire n_1123;
wire n_1122;
wire n_768;
wire n_1125;
wire n_1124;
wire n_1127;
wire n_1126;
wire n_1129;
wire n_1128;
wire n_1077;
wire n_1131;
wire n_1130;
wire n_1133;
wire n_1132;
wire n_1135;
wire n_1134;
wire n_1137;
wire n_1136;
wire n_2197;
wire n_2226;
wire n_2256;
wire n_1139;
wire n_1138;
wire n_2284;
wire n_2313;
wire n_2343;
wire n_1141;
wire n_1140;
wire n_2371;
wire n_2400;
wire n_2430;
wire n_1143;
wire n_1142;
wire n_2458;
wire n_2487;
wire n_2517;
wire n_1145;
wire n_1144;
wire n_2545;
wire n_2574;
wire n_2604;
wire n_1147;
wire n_1146;
wire n_2632;
wire n_2661;
wire n_2691;
wire n_1149;
wire n_1148;
wire n_2719;
wire n_2748;
wire n_2778;
wire n_1151;
wire n_1150;
wire n_1153;
wire n_1152;
wire n_1155;
wire n_1154;
wire n_2107;
wire n_1157;
wire n_1156;
wire n_2100;
wire n_1159;
wire n_1158;
wire n_2085;
wire n_1161;
wire n_1160;
wire n_1163;
wire n_1162;
wire n_2094;
wire n_1165;
wire n_1164;
wire n_1167;
wire n_1166;
wire n_1169;
wire n_1168;
wire n_1171;
wire n_1170;
wire n_1173;
wire n_1172;
wire n_1175;
wire n_1174;
wire n_1177;
wire n_1176;
wire n_1179;
wire n_1178;
wire n_1181;
wire n_1180;
wire n_1183;
wire n_1182;
wire n_1185;
wire n_1184;
wire n_2196;
wire n_2225;
wire n_2255;
wire n_1187;
wire n_1186;
wire n_2283;
wire n_2312;
wire n_2342;
wire n_1189;
wire n_1188;
wire n_2370;
wire n_2399;
wire n_2429;
wire n_1191;
wire n_1190;
wire n_2457;
wire n_2486;
wire n_2516;
wire n_1193;
wire n_1192;
wire n_2544;
wire n_2573;
wire n_2603;
wire n_1195;
wire n_1194;
wire n_2631;
wire n_2660;
wire n_2690;
wire n_1197;
wire n_1196;
wire n_2718;
wire n_2747;
wire n_2777;
wire n_1199;
wire n_1198;
wire n_1201;
wire n_1200;
wire n_1203;
wire n_1202;
wire n_2092;
wire n_1205;
wire n_1204;
wire n_2071;
wire n_1207;
wire n_1206;
wire n_1209;
wire n_1208;
wire n_1211;
wire n_1210;
wire n_2079;
wire n_1213;
wire n_1212;
wire n_1215;
wire n_1214;
wire n_1217;
wire n_1216;
wire n_1219;
wire n_1218;
wire n_1221;
wire n_1220;
wire n_1223;
wire n_1222;
wire n_1225;
wire n_1224;
wire n_1227;
wire n_1226;
wire n_1229;
wire n_1228;
wire n_1231;
wire n_1230;
wire n_2195;
wire n_2224;
wire n_2254;
wire n_1233;
wire n_1232;
wire n_2282;
wire n_2311;
wire n_2341;
wire n_1235;
wire n_1234;
wire n_2369;
wire n_2398;
wire n_2428;
wire n_1237;
wire n_1236;
wire n_2456;
wire n_2485;
wire n_2515;
wire n_1239;
wire n_1238;
wire n_2543;
wire n_2572;
wire n_2602;
wire n_1241;
wire n_1240;
wire n_2630;
wire n_2659;
wire n_2689;
wire n_1243;
wire n_1242;
wire n_2717;
wire n_2746;
wire n_2776;
wire n_1245;
wire n_1244;
wire n_1247;
wire n_1246;
wire n_2077;
wire n_1249;
wire n_1248;
wire n_2070;
wire n_1251;
wire n_1250;
wire n_1253;
wire n_1252;
wire n_1255;
wire n_1254;
wire n_2064;
wire n_1257;
wire n_1256;
wire n_2057;
wire n_1259;
wire n_1258;
wire n_1261;
wire n_1260;
wire n_1263;
wire n_1262;
wire n_1265;
wire n_1264;
wire n_1267;
wire n_1266;
wire n_1269;
wire n_1268;
wire n_1271;
wire n_1270;
wire n_1273;
wire n_1272;
wire n_1275;
wire n_1274;
wire n_2194;
wire n_2223;
wire n_2253;
wire n_1277;
wire n_1276;
wire n_2281;
wire n_2310;
wire n_2340;
wire n_1279;
wire n_1278;
wire n_2368;
wire n_2397;
wire n_2427;
wire n_1281;
wire n_1280;
wire n_2455;
wire n_2484;
wire n_2514;
wire n_1283;
wire n_1282;
wire n_2542;
wire n_2571;
wire n_2601;
wire n_1285;
wire n_1284;
wire n_2629;
wire n_2658;
wire n_2688;
wire n_1287;
wire n_1286;
wire n_1289;
wire n_1288;
wire n_1291;
wire n_1290;
wire n_2062;
wire n_1293;
wire n_1292;
wire n_2055;
wire n_2040;
wire n_1295;
wire n_1294;
wire n_1297;
wire n_1296;
wire n_1299;
wire n_1298;
wire n_2049;
wire n_1301;
wire n_1300;
wire n_1303;
wire n_1302;
wire n_1305;
wire n_1304;
wire n_1307;
wire n_1306;
wire n_1309;
wire n_1308;
wire n_1311;
wire n_1310;
wire n_1313;
wire n_1312;
wire n_1315;
wire n_1314;
wire n_1317;
wire n_1316;
wire n_2193;
wire n_2222;
wire n_2252;
wire n_1319;
wire n_1318;
wire n_2280;
wire n_2309;
wire n_2339;
wire n_1321;
wire n_1320;
wire n_2367;
wire n_2396;
wire n_2426;
wire n_1323;
wire n_1322;
wire n_2454;
wire n_2483;
wire n_2513;
wire n_1325;
wire n_1324;
wire n_2541;
wire n_2570;
wire n_2600;
wire n_1327;
wire n_1326;
wire n_2628;
wire n_2657;
wire n_2687;
wire n_1329;
wire n_1328;
wire n_1331;
wire n_1330;
wire n_1333;
wire n_1332;
wire n_2047;
wire n_1335;
wire n_1334;
wire n_2027;
wire n_1337;
wire n_1336;
wire n_1339;
wire n_1338;
wire n_2034;
wire n_1341;
wire n_1340;
wire n_1343;
wire n_1342;
wire n_1345;
wire n_1344;
wire n_1347;
wire n_1346;
wire n_1349;
wire n_1348;
wire n_1351;
wire n_1350;
wire n_1353;
wire n_1352;
wire n_1355;
wire n_1354;
wire n_1357;
wire n_1356;
wire n_2192;
wire n_2221;
wire n_2251;
wire n_1359;
wire n_1358;
wire n_2279;
wire n_2308;
wire n_2338;
wire n_1361;
wire n_1360;
wire n_2366;
wire n_2395;
wire n_2425;
wire n_1363;
wire n_1362;
wire n_2453;
wire n_2482;
wire n_2512;
wire n_1365;
wire n_1364;
wire n_2540;
wire n_2569;
wire n_2599;
wire n_1367;
wire n_1366;
wire n_2627;
wire n_2656;
wire n_2686;
wire n_1369;
wire n_1368;
wire n_1371;
wire n_1370;
wire n_2032;
wire n_1373;
wire n_1372;
wire n_2025;
wire n_1375;
wire n_1374;
wire n_1377;
wire n_1376;
wire n_2019;
wire n_1379;
wire n_1378;
wire n_1381;
wire n_1380;
wire n_2012;
wire n_1383;
wire n_1382;
wire n_1385;
wire n_1384;
wire n_1387;
wire n_1386;
wire n_1389;
wire n_1388;
wire n_1391;
wire n_1390;
wire n_1393;
wire n_1392;
wire n_1395;
wire n_1394;
wire n_2191;
wire n_2220;
wire n_2250;
wire n_1397;
wire n_1396;
wire n_2278;
wire n_2307;
wire n_2337;
wire n_1399;
wire n_1398;
wire n_2365;
wire n_2394;
wire n_2424;
wire n_1401;
wire n_1400;
wire n_2452;
wire n_2481;
wire n_2511;
wire n_1403;
wire n_1402;
wire n_2539;
wire n_2568;
wire n_2598;
wire n_1405;
wire n_1404;
wire n_1407;
wire n_1406;
wire n_1409;
wire n_1408;
wire n_2017;
wire n_2010;
wire n_1411;
wire n_1410;
wire n_1995;
wire n_1413;
wire n_1412;
wire n_1415;
wire n_1414;
wire n_2004;
wire n_1417;
wire n_1416;
wire n_1419;
wire n_1418;
wire n_1421;
wire n_1420;
wire n_1423;
wire n_1422;
wire n_1425;
wire n_1424;
wire n_1427;
wire n_1426;
wire n_1429;
wire n_1428;
wire n_1431;
wire n_1430;
wire n_2190;
wire n_2219;
wire n_2249;
wire n_1433;
wire n_1432;
wire n_2277;
wire n_2306;
wire n_2336;
wire n_1435;
wire n_1434;
wire n_2364;
wire n_2393;
wire n_2423;
wire n_1437;
wire n_1436;
wire n_2451;
wire n_2480;
wire n_2510;
wire n_1439;
wire n_1438;
wire n_2538;
wire n_2567;
wire n_2597;
wire n_1441;
wire n_1440;
wire n_1443;
wire n_1442;
wire n_2002;
wire n_1445;
wire n_1444;
wire n_1981;
wire n_1447;
wire n_1446;
wire n_1449;
wire n_1448;
wire n_1989;
wire n_1451;
wire n_1450;
wire n_1453;
wire n_1452;
wire n_1455;
wire n_1454;
wire n_1457;
wire n_1456;
wire n_1459;
wire n_1458;
wire n_1461;
wire n_1460;
wire n_1463;
wire n_1462;
wire n_1465;
wire n_1464;
wire n_2189;
wire n_2218;
wire n_2248;
wire n_1467;
wire n_1466;
wire n_2276;
wire n_2305;
wire n_2335;
wire n_1469;
wire n_1468;
wire n_2363;
wire n_2392;
wire n_2422;
wire n_1471;
wire n_1470;
wire n_2450;
wire n_2479;
wire n_2509;
wire n_1473;
wire n_1472;
wire n_2537;
wire n_2566;
wire n_2596;
wire n_1475;
wire n_1474;
wire n_1477;
wire n_1476;
wire n_1987;
wire n_1479;
wire n_1478;
wire n_1980;
wire n_1481;
wire n_1480;
wire n_1483;
wire n_1482;
wire n_1974;
wire n_1967;
wire n_1485;
wire n_1484;
wire n_1487;
wire n_1486;
wire n_1489;
wire n_1488;
wire n_1491;
wire n_1490;
wire n_1493;
wire n_1492;
wire n_1495;
wire n_1494;
wire n_1497;
wire n_1496;
wire n_2188;
wire n_2217;
wire n_2247;
wire n_1499;
wire n_1498;
wire n_2275;
wire n_2304;
wire n_2334;
wire n_1501;
wire n_1500;
wire n_2362;
wire n_2391;
wire n_2421;
wire n_1503;
wire n_1502;
wire n_2449;
wire n_2478;
wire n_2508;
wire n_1505;
wire n_1504;
wire n_1507;
wire n_1506;
wire n_1972;
wire n_1509;
wire n_1508;
wire n_1965;
wire n_1950;
wire n_1511;
wire n_1510;
wire n_1513;
wire n_1512;
wire n_1959;
wire n_1515;
wire n_1514;
wire n_1517;
wire n_1516;
wire n_1519;
wire n_1518;
wire n_1521;
wire n_1520;
wire n_1523;
wire n_1522;
wire n_1525;
wire n_1524;
wire n_1527;
wire n_1526;
wire n_2187;
wire n_2216;
wire n_2246;
wire n_1529;
wire n_1528;
wire n_2274;
wire n_2303;
wire n_2333;
wire n_1531;
wire n_1530;
wire n_2361;
wire n_2390;
wire n_2420;
wire n_1533;
wire n_1532;
wire n_2448;
wire n_2477;
wire n_2507;
wire n_1535;
wire n_1534;
wire n_1537;
wire n_1536;
wire n_1957;
wire n_1539;
wire n_1538;
wire n_1937;
wire n_1541;
wire n_1540;
wire n_1543;
wire n_1542;
wire n_1944;
wire n_1545;
wire n_1544;
wire n_1547;
wire n_1546;
wire n_1549;
wire n_1548;
wire n_1551;
wire n_1550;
wire n_1553;
wire n_1552;
wire n_1555;
wire n_1554;
wire n_2186;
wire n_2215;
wire n_2245;
wire n_1557;
wire n_1556;
wire n_2273;
wire n_2302;
wire n_2332;
wire n_1559;
wire n_1558;
wire n_2360;
wire n_2389;
wire n_2419;
wire n_1561;
wire n_1560;
wire n_2447;
wire n_2476;
wire n_2506;
wire n_1563;
wire n_1562;
wire n_1942;
wire n_1565;
wire n_1564;
wire n_1935;
wire n_1567;
wire n_1566;
wire n_1569;
wire n_1568;
wire n_1929;
wire n_1571;
wire n_1570;
wire n_1922;
wire n_1573;
wire n_1572;
wire n_1575;
wire n_1574;
wire n_1577;
wire n_1576;
wire n_1579;
wire n_1578;
wire n_1581;
wire n_1580;
wire n_2185;
wire n_2214;
wire n_2244;
wire n_1583;
wire n_1582;
wire n_2272;
wire n_2301;
wire n_2331;
wire n_1585;
wire n_1584;
wire n_2359;
wire n_2388;
wire n_2418;
wire n_1587;
wire n_1586;
wire n_1589;
wire n_1588;
wire n_1927;
wire n_1591;
wire n_1590;
wire n_1920;
wire n_1905;
wire n_1593;
wire n_1592;
wire n_1914;
wire n_1595;
wire n_1594;
wire n_1597;
wire n_1596;
wire n_1599;
wire n_1598;
wire n_1601;
wire n_1600;
wire n_1603;
wire n_1602;
wire n_1605;
wire n_1604;
wire n_2184;
wire n_2213;
wire n_2243;
wire n_1607;
wire n_1606;
wire n_2271;
wire n_2300;
wire n_2330;
wire n_1609;
wire n_1608;
wire n_2358;
wire n_2387;
wire n_2417;
wire n_1611;
wire n_1610;
wire n_1613;
wire n_1612;
wire n_1912;
wire n_1892;
wire n_1615;
wire n_1614;
wire n_1617;
wire n_1616;
wire n_1899;
wire n_1619;
wire n_1618;
wire n_1621;
wire n_1620;
wire n_1623;
wire n_1622;
wire n_1625;
wire n_1624;
wire n_1627;
wire n_1626;
wire n_2183;
wire n_2212;
wire n_2242;
wire n_1629;
wire n_1628;
wire n_2270;
wire n_2299;
wire n_2329;
wire n_1631;
wire n_1630;
wire n_2357;
wire n_2386;
wire n_2416;
wire n_1633;
wire n_1632;
wire n_1897;
wire n_1635;
wire n_1634;
wire n_1890;
wire n_1637;
wire n_1636;
wire n_1884;
wire n_1639;
wire n_1638;
wire n_1877;
wire n_1641;
wire n_1640;
wire n_1643;
wire n_1642;
wire n_1645;
wire n_1644;
wire n_1647;
wire n_1646;
wire n_2182;
wire n_2211;
wire n_2241;
wire n_1649;
wire n_1648;
wire n_2269;
wire n_2298;
wire n_2328;
wire n_1651;
wire n_1650;
wire n_1653;
wire n_1652;
wire n_1882;
wire n_1875;
wire n_1860;
wire n_1655;
wire n_1654;
wire n_1869;
wire n_1657;
wire n_1656;
wire n_1659;
wire n_1658;
wire n_1661;
wire n_1660;
wire n_1663;
wire n_1662;
wire n_1665;
wire n_1664;
wire n_2181;
wire n_2210;
wire n_2240;
wire n_1667;
wire n_1666;
wire n_2268;
wire n_2297;
wire n_2327;
wire n_1669;
wire n_1668;
wire n_1867;
wire n_1671;
wire n_1670;
wire n_1846;
wire n_1673;
wire n_1672;
wire n_1854;
wire n_1675;
wire n_1674;
wire n_1677;
wire n_1676;
wire n_1679;
wire n_1678;
wire n_1681;
wire n_1680;
wire n_2180;
wire n_2209;
wire n_2239;
wire n_1683;
wire n_1682;
wire n_2267;
wire n_2296;
wire n_2326;
wire n_1685;
wire n_1684;
wire n_1852;
wire n_1845;
wire n_1687;
wire n_1686;
wire n_1839;
wire n_1689;
wire n_1688;
wire n_1832;
wire n_1691;
wire n_1690;
wire n_1693;
wire n_1692;
wire n_1695;
wire n_1694;
wire n_2179;
wire n_2208;
wire n_2238;
wire n_1697;
wire n_1696;
wire n_1837;
wire n_1699;
wire n_1698;
wire n_1830;
wire n_1815;
wire n_1701;
wire n_1700;
wire n_1824;
wire n_1703;
wire n_1702;
wire n_1705;
wire n_1704;
wire n_1707;
wire n_1706;
wire n_2178;
wire n_2207;
wire n_2237;
wire n_1709;
wire n_1708;
wire n_1822;
wire n_1711;
wire n_1710;
wire n_1803;
wire n_1808;
wire n_1713;
wire n_1712;
wire n_1715;
wire n_1714;
wire n_1717;
wire n_1716;
wire n_2177;
wire n_2206;
wire n_2236;
wire n_1719;
wire n_1718;
wire n_1801;
wire n_1795;
wire n_1721;
wire n_1720;
wire n_1787;
wire n_1723;
wire n_1722;
wire n_1725;
wire n_1724;
wire n_1793;
wire n_1786;
wire n_1727;
wire n_1726;
wire n_1771;
wire n_1780;
wire n_1729;
wire n_1728;
wire n_1731;
wire n_1730;
wire n_1778;
wire n_1758;
wire n_1764;
wire n_1733;
wire n_1732;
wire n_1735;
wire n_1734;
wire n_1752;
wire n_1743;
wire n_1737;
wire n_1736;
wire n_1745;
wire n_3464;
wire n_3470;
wire n_3481;
wire n_3471;
wire n_3482;
wire n_1753;
wire n_3483;
wire n_3485;
wire n_3484;
wire n_1760;
wire n_3472;
wire n_3478;
wire n_3480;
wire n_3479;
wire n_3467;
wire n_1765;
wire n_3466;
wire n_3469;
wire n_3468;
wire n_1774;
wire n_3474;
wire n_3476;
wire n_3475;
wire n_1782;
wire n_1779;
wire n_1785;
wire n_1784;
wire n_1783;
wire n_1781;
wire n_3444;
wire n_2172;
wire n_3443;
wire n_3404;
wire n_1791;
wire n_1790;
wire n_1788;
wire n_1789;
wire n_1813;
wire n_1812;
wire n_1814;
wire n_1810;
wire n_1792;
wire n_1797;
wire n_1794;
wire n_1800;
wire n_1799;
wire n_1798;
wire n_1796;
wire n_2171;
wire n_1802;
wire n_1821;
wire n_1807;
wire n_1806;
wire n_1804;
wire n_1805;
wire n_1819;
wire n_1818;
wire n_1816;
wire n_3438;
wire n_3410;
wire n_1809;
wire n_1811;
wire n_2170;
wire n_1817;
wire n_3437;
wire n_1820;
wire n_3405;
wire n_1826;
wire n_1823;
wire n_1829;
wire n_1828;
wire n_1827;
wire n_1825;
wire n_2169;
wire n_1834;
wire n_1831;
wire n_1835;
wire n_1833;
wire n_1836;
wire n_1841;
wire n_1838;
wire n_1844;
wire n_1843;
wire n_1842;
wire n_1840;
wire n_2166;
wire n_1866;
wire n_1851;
wire n_1849;
wire n_1847;
wire n_1848;
wire n_1865;
wire n_1861;
wire n_1850;
wire n_3435;
wire n_1856;
wire n_1853;
wire n_1859;
wire n_1858;
wire n_1857;
wire n_1855;
wire n_2164;
wire n_1863;
wire n_1862;
wire n_1864;
wire n_3434;
wire n_1871;
wire n_1868;
wire n_1874;
wire n_1873;
wire n_1872;
wire n_1870;
wire n_2163;
wire n_1879;
wire n_1876;
wire n_1880;
wire n_1878;
wire n_1881;
wire n_1886;
wire n_1883;
wire n_1889;
wire n_1888;
wire n_1887;
wire n_1885;
wire n_2162;
wire n_1891;
wire n_1911;
wire n_1896;
wire n_1895;
wire n_1893;
wire n_1894;
wire n_1909;
wire n_1908;
wire n_1906;
wire n_3432;
wire n_1901;
wire n_1898;
wire n_1904;
wire n_1903;
wire n_1902;
wire n_1900;
wire n_2158;
wire n_1907;
wire n_3431;
wire n_1910;
wire n_1916;
wire n_1913;
wire n_1919;
wire n_1918;
wire n_1917;
wire n_1915;
wire n_2156;
wire n_1924;
wire n_1921;
wire n_1925;
wire n_1923;
wire n_1926;
wire n_1931;
wire n_1928;
wire n_1934;
wire n_1933;
wire n_1932;
wire n_1930;
wire n_2155;
wire n_1936;
wire n_1956;
wire n_1941;
wire n_1940;
wire n_1938;
wire n_1939;
wire n_1954;
wire n_1953;
wire n_1951;
wire n_3429;
wire n_1946;
wire n_1943;
wire n_1949;
wire n_1948;
wire n_1947;
wire n_1945;
wire n_2154;
wire n_1952;
wire n_3428;
wire n_1955;
wire n_1961;
wire n_1958;
wire n_1964;
wire n_1963;
wire n_1962;
wire n_1960;
wire n_2152;
wire n_1969;
wire n_1966;
wire n_1970;
wire n_1968;
wire n_1971;
wire n_1976;
wire n_1973;
wire n_1979;
wire n_1978;
wire n_1977;
wire n_1975;
wire n_2151;
wire n_2001;
wire n_1986;
wire n_1984;
wire n_1982;
wire n_1983;
wire n_2000;
wire n_1996;
wire n_1985;
wire n_3426;
wire n_1991;
wire n_1988;
wire n_1994;
wire n_1993;
wire n_1992;
wire n_1990;
wire n_2150;
wire n_1998;
wire n_1997;
wire n_1999;
wire n_3422;
wire n_2006;
wire n_2003;
wire n_2009;
wire n_2008;
wire n_2007;
wire n_2005;
wire n_2149;
wire n_2014;
wire n_2011;
wire n_2015;
wire n_2013;
wire n_2016;
wire n_2021;
wire n_2018;
wire n_2024;
wire n_2023;
wire n_2022;
wire n_2020;
wire n_2148;
wire n_2026;
wire n_2046;
wire n_2031;
wire n_2030;
wire n_2028;
wire n_2029;
wire n_2044;
wire n_2043;
wire n_2041;
wire n_3420;
wire n_2036;
wire n_2033;
wire n_2039;
wire n_2038;
wire n_2037;
wire n_2035;
wire n_2146;
wire n_2042;
wire n_3419;
wire n_2045;
wire n_2051;
wire n_2048;
wire n_2054;
wire n_2053;
wire n_2052;
wire n_2050;
wire n_2144;
wire n_2059;
wire n_2056;
wire n_2060;
wire n_2058;
wire n_2061;
wire n_2066;
wire n_2063;
wire n_2069;
wire n_2068;
wire n_2067;
wire n_2065;
wire n_2143;
wire n_2091;
wire n_2076;
wire n_2074;
wire n_2072;
wire n_2073;
wire n_2090;
wire n_2086;
wire n_2075;
wire n_3417;
wire n_2081;
wire n_2078;
wire n_2084;
wire n_2083;
wire n_2082;
wire n_2080;
wire n_2142;
wire n_2088;
wire n_2087;
wire n_2089;
wire n_3416;
wire n_2096;
wire n_2093;
wire n_2099;
wire n_2098;
wire n_2097;
wire n_2095;
wire n_2141;
wire n_2104;
wire n_2101;
wire n_2105;
wire n_2103;
wire n_2106;
wire n_2111;
wire n_2108;
wire n_2114;
wire n_2113;
wire n_2112;
wire n_2110;
wire n_2138;
wire n_1762;
wire n_2121;
wire n_2119;
wire n_2117;
wire n_2118;
wire n_1761;
wire n_2131;
wire n_2120;
wire n_3414;
wire n_2127;
wire n_2123;
wire n_2132;
wire n_2129;
wire n_2128;
wire n_1759;
wire n_1757;
wire n_1767;
wire n_2140;
wire n_1768;
wire n_1770;
wire n_1769;
wire n_1777;
wire n_2126;
wire n_2125;
wire n_984;
wire n_2160;
wire n_1763;
wire n_2161;
wire n_1766;
wire n_1772;
wire n_2168;
wire n_1773;
wire n_1776;
wire n_1775;
wire n_3425;
wire n_2135;
wire n_2133;
wire n_3442;
wire n_2136;
wire n_2134;
wire n_3441;
wire n_3440;
wire n_3406;
wire n_3439;
wire n_3436;
wire n_3433;
wire n_3430;
wire n_3427;
wire n_3421;
wire n_3418;
wire n_3415;
wire n_3413;
wire n_3412;
wire n_3411;
wire n_3042;
wire n_3396;
wire n_3399;
wire n_3398;
wire n_3043;
wire n_3395;
wire n_3401;
wire n_3394;
wire n_3044;
wire n_3402;
wire n_3392;
wire n_3045;
wire n_3391;
wire n_3052;
wire n_3051;
wire n_3048;
wire n_3049;
wire n_3046;
wire n_3388;
wire n_3379;
wire n_3053;
wire n_3047;
wire n_3389;
wire n_3383;
wire n_3050;
wire n_3386;
wire n_3384;
wire n_3390;
wire n_3381;
wire n_3377;
wire n_3060;
wire n_3059;
wire n_3056;
wire n_3057;
wire n_3054;
wire n_3374;
wire n_3365;
wire n_3061;
wire n_3055;
wire n_3375;
wire n_3369;
wire n_3058;
wire n_3372;
wire n_3370;
wire n_3376;
wire n_3367;
wire n_3363;
wire n_3068;
wire n_3067;
wire n_3064;
wire n_3065;
wire n_3062;
wire n_3360;
wire n_3351;
wire n_3069;
wire n_3063;
wire n_3361;
wire n_3355;
wire n_3066;
wire n_3358;
wire n_3356;
wire n_3362;
wire n_3353;
wire n_3349;
wire n_3076;
wire n_3075;
wire n_3072;
wire n_3073;
wire n_3070;
wire n_3315;
wire n_3305;
wire n_3077;
wire n_3071;
wire n_3314;
wire n_3317;
wire n_3307;
wire n_3074;
wire n_3316;
wire n_3312;
wire n_3309;
wire n_3319;
wire n_3105;
wire n_3084;
wire n_3083;
wire n_3080;
wire n_3081;
wire n_3078;
wire n_3343;
wire n_3287;
wire n_3085;
wire n_3079;
wire n_3342;
wire n_3345;
wire n_3289;
wire n_3082;
wire n_3344;
wire n_3348;
wire n_3291;
wire n_3347;
wire n_3103;
wire n_3092;
wire n_3091;
wire n_3088;
wire n_3089;
wire n_3086;
wire n_3326;
wire n_3299;
wire n_3093;
wire n_3087;
wire n_3325;
wire n_3328;
wire n_3301;
wire n_3090;
wire n_3327;
wire n_3323;
wire n_3303;
wire n_3330;
wire n_3101;
wire n_3100;
wire n_3099;
wire n_3096;
wire n_3097;
wire n_3094;
wire n_3335;
wire n_3293;
wire n_3107;
wire n_3095;
wire n_3334;
wire n_3337;
wire n_3296;
wire n_3098;
wire n_3336;
wire n_3332;
wire n_3297;
wire n_3102;
wire n_3298;
wire n_3322;
wire n_3104;
wire n_3286;
wire n_3340;
wire n_3106;
wire n_3304;
wire n_3311;
wire n_3338;
wire n_3424;
wire n_3423;
wire n_3284;
wire n_3114;
wire n_3113;
wire n_3110;
wire n_3111;
wire n_3108;
wire n_3253;
wire n_3243;
wire n_3115;
wire n_3109;
wire n_3252;
wire n_3255;
wire n_3245;
wire n_3112;
wire n_3254;
wire n_3250;
wire n_3247;
wire n_3257;
wire n_3143;
wire n_3122;
wire n_3121;
wire n_3118;
wire n_3119;
wire n_3116;
wire n_3278;
wire n_3236;
wire n_3123;
wire n_3117;
wire n_3277;
wire n_3280;
wire n_3238;
wire n_3120;
wire n_3279;
wire n_3283;
wire n_3240;
wire n_3282;
wire n_3141;
wire n_3130;
wire n_3129;
wire n_3126;
wire n_3127;
wire n_3124;
wire n_3264;
wire n_3222;
wire n_3131;
wire n_3125;
wire n_3263;
wire n_3266;
wire n_3224;
wire n_3128;
wire n_3265;
wire n_3261;
wire n_3226;
wire n_3268;
wire n_3140;
wire n_3139;
wire n_3137;
wire n_3136;
wire n_3133;
wire n_3132;
wire n_3232;
wire n_3272;
wire n_3229;
wire n_3145;
wire n_3134;
wire n_3135;
wire n_3271;
wire n_3230;
wire n_3138;
wire n_3273;
wire n_3233;
wire n_3234;
wire n_3221;
wire n_3260;
wire n_3142;
wire n_3235;
wire n_3275;
wire n_3144;
wire n_3242;
wire n_3249;
wire n_3274;
wire n_3219;
wire n_3152;
wire n_3151;
wire n_3148;
wire n_3149;
wire n_3146;
wire n_3216;
wire n_3207;
wire n_3153;
wire n_3147;
wire n_3217;
wire n_3211;
wire n_3150;
wire n_3214;
wire n_3212;
wire n_3218;
wire n_3209;
wire n_3205;
wire n_3160;
wire n_3159;
wire n_3156;
wire n_3157;
wire n_3154;
wire n_3202;
wire n_3193;
wire n_3161;
wire n_3155;
wire n_3203;
wire n_3197;
wire n_3158;
wire n_3200;
wire n_3198;
wire n_3204;
wire n_3195;
wire n_3191;
wire n_3169;
wire n_3168;
wire n_3167;
wire n_3163;
wire n_3162;
wire n_3181;
wire n_3188;
wire n_3170;
wire n_3164;
wire n_3165;
wire n_3166;
wire n_3177;
wire n_3189;
wire n_3185;
wire n_3183;
wire n_3182;
wire n_3190;
wire n_3178;
wire n_3175;
wire n_3171;
wire n_3450;
wire n_3486;
wire n_3451;
wire n_3173;
wire n_3172;
wire n_3407;
wire n_3454;
wire n_3408;
wire n_3455;
wire n_3409;
wire n_3174;
wire n_3176;
wire n_3179;
wire n_3184;
wire n_3446;
wire n_3180;
wire n_3187;
wire n_3186;
wire n_3192;
wire n_3196;
wire n_3199;
wire n_3194;
wire n_3201;
wire n_3206;
wire n_3210;
wire n_3213;
wire n_3208;
wire n_3215;
wire n_3241;
wire n_3220;
wire n_3248;
wire n_3227;
wire n_3269;
wire n_3259;
wire n_3223;
wire n_3267;
wire n_3262;
wire n_3225;
wire n_3228;
wire n_3231;
wire n_3270;
wire n_3237;
wire n_3281;
wire n_3276;
wire n_3239;
wire n_3258;
wire n_3244;
wire n_3256;
wire n_3251;
wire n_3246;
wire n_3292;
wire n_3285;
wire n_3310;
wire n_3320;
wire n_3321;
wire n_3331;
wire n_3288;
wire n_3346;
wire n_3341;
wire n_3290;
wire n_3333;
wire n_3295;
wire n_3339;
wire n_3294;
wire n_3300;
wire n_3329;
wire n_3324;
wire n_3302;
wire n_3306;
wire n_3318;
wire n_3313;
wire n_3308;
wire n_3350;
wire n_3354;
wire n_3357;
wire n_3352;
wire n_3359;
wire n_3364;
wire n_3368;
wire n_3371;
wire n_3366;
wire n_3373;
wire n_3378;
wire n_3382;
wire n_3385;
wire n_3380;
wire n_3387;
wire n_3403;
wire n_3393;
wire n_3400;
wire n_3456;
wire n_3453;
wire n_3457;
wire n_2289;
wire n_2318;
wire n_2348;
wire n_873;
wire n_872;
wire n_2202;
wire n_2231;
wire n_2261;
wire n_871;
wire n_2165;
wire n_949;
wire n_948;
wire n_2550;
wire n_2579;
wire n_2609;
wire n_879;
wire n_878;
wire n_2463;
wire n_2492;
wire n_2522;
wire n_877;
wire n_876;
wire n_2376;
wire n_2405;
wire n_2435;
wire n_875;
wire n_874;
wire n_947;
wire n_946;
wire n_1005;
wire n_1004;
wire n_2287;
wire n_2316;
wire n_2346;
wire n_985;
wire n_2200;
wire n_2229;
wire n_2259;
wire n_983;
wire n_2137;
wire n_1056;
wire n_2124;
wire n_1066;
wire n_2811;
wire n_2840;
wire n_2870;
wire n_885;
wire n_2724;
wire n_2753;
wire n_2783;
wire n_883;
wire n_882;
wire n_2637;
wire n_2666;
wire n_2696;
wire n_881;
wire n_880;
wire n_945;
wire n_944;
wire n_901;
wire n_899;
wire n_963;
wire n_2524;
wire n_2552;
wire n_2581;
wire n_765;
wire n_2437;
wire n_2465;
wire n_2494;
wire n_763;
wire n_2350;
wire n_2378;
wire n_2407;
wire n_761;
wire n_837;
wire n_2785;
wire n_2813;
wire n_2842;
wire n_771;
wire n_2698;
wire n_2726;
wire n_2755;
wire n_769;
wire n_2611;
wire n_2639;
wire n_2668;
wire n_767;
wire n_835;
wire n_2958;
wire n_2987;
wire n_3015;
wire n_775;
wire n_2872;
wire n_2900;
wire n_2929;
wire n_773;
wire n_3014;
wire n_833;
wire n_895;
wire n_961;
wire n_1021;
wire n_2782;
wire n_2810;
wire n_2839;
wire n_940;
wire n_2695;
wire n_2723;
wire n_2752;
wire n_938;
wire n_2608;
wire n_2636;
wire n_2665;
wire n_936;
wire n_955;
wire n_2928;
wire n_2957;
wire n_2986;
wire n_2898;
wire n_2927;
wire n_2956;
wire n_887;
wire n_2869;
wire n_2897;
wire n_2926;
wire n_942;
wire n_2157;
wire n_2147;
wire n_953;
wire n_2145;
wire n_2130;
wire n_1006;
wire n_1019;
wire n_1738;
wire n_1741;
wire n_1747;
wire n_1748;
wire n_1744;
wire n_1746;
wire n_1749;
wire n_1751;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_3445;
wire n_1750;
wire n_1740;
wire n_1742;
wire n_1739;
wire n_3447;
wire n_3458;
wire n_3448;
wire n_3461;
wire n_3460;
wire n_3449;
wire n_3452;
wire n_3462;
wire n_3459;
wire n_3463;
wire n_3465;
wire n_3477;
wire n_3473;


INV_X1 i_2680 (.ZN (n_3486), .A (n_1739));
NAND2_X1 i_2679 (.ZN (n_3485), .A1 (inputB[31]), .A2 (inputA[28]));
NOR2_X1 i_2678 (.ZN (n_3484), .A1 (n_3444), .A2 (n_3405));
NAND2_X1 i_2677 (.ZN (n_3483), .A1 (n_3485), .A2 (n_3484));
NOR2_X1 i_2676 (.ZN (n_3482), .A1 (n_3443), .A2 (n_3406));
NAND2_X1 i_2675 (.ZN (n_3481), .A1 (inputB[28]), .A2 (inputA[31]));
NAND2_X1 i_2674 (.ZN (n_3480), .A1 (inputB[28]), .A2 (inputA[30]));
NOR2_X1 i_2673 (.ZN (n_3479), .A1 (n_3410), .A2 (n_3441));
NAND2_X1 i_2672 (.ZN (n_3478), .A1 (n_3480), .A2 (n_3479));
INV_X1 i_2671 (.ZN (n_3477), .A (n_3478));
NOR3_X1 i_2670 (.ZN (n_3476), .A1 (n_3441), .A2 (n_3480), .A3 (n_3405));
AOI22_X1 i_2669 (.ZN (n_3475), .A1 (inputB[28]), .A2 (inputA[29]), .B1 (inputB[27]), .B2 (inputA[30]));
NOR2_X1 i_2668 (.ZN (n_3474), .A1 (n_3410), .A2 (n_3440));
NOR2_X1 i_2667 (.ZN (n_3473), .A1 (n_3475), .A2 (n_3474));
NOR2_X1 i_2666 (.ZN (n_3472), .A1 (n_3476), .A2 (n_3473));
OAI22_X1 i_2665 (.ZN (n_3471), .A1 (n_3480), .A2 (n_3479), .B1 (n_3477), .B2 (n_3472));
NOR2_X1 i_2664 (.ZN (n_3470), .A1 (n_3481), .A2 (n_3471));
NAND2_X1 i_2663 (.ZN (n_3469), .A1 (inputB[31]), .A2 (inputA[27]));
NOR2_X1 i_2662 (.ZN (n_3468), .A1 (n_3444), .A2 (n_3404));
NOR2_X1 i_2661 (.ZN (n_3467), .A1 (n_3405), .A2 (n_3443));
NAND2_X1 i_2660 (.ZN (n_3466), .A1 (n_3469), .A2 (n_3468));
INV_X1 i_2659 (.ZN (n_3465), .A (n_3466));
OAI22_X1 i_2658 (.ZN (n_3464), .A1 (n_3469), .A2 (n_3468), .B1 (n_3467), .B2 (n_3465));
NOR2_X1 i_2657 (.ZN (n_3463), .A1 (n_3444), .A2 (n_3406));
INV_X1 i_2656 (.ZN (n_3462), .A (n_3463));
AOI21_X1 i_2655 (.ZN (n_3461), .A (n_3462), .B1 (inputB[29]), .B2 (inputA[31]));
NOR3_X1 i_2654 (.ZN (n_3460), .A1 (n_3443), .A2 (n_3463), .A3 (n_3410));
INV_X1 i_2653 (.ZN (n_3459), .A (n_3460));
NAND2_X1 i_2652 (.ZN (n_3458), .A1 (inputB[31]), .A2 (inputA[29]));
AOI21_X1 i_2651 (.ZN (n_3457), .A (n_3461), .B1 (n_3459), .B2 (n_3458));
OAI22_X1 i_2650 (.ZN (n_3456), .A1 (n_3406), .A2 (n_3445), .B1 (n_3444), .B2 (n_3410));
NOR2_X1 i_2649 (.ZN (n_3455), .A1 (n_3410), .A2 (n_3445));
INV_X1 i_2648 (.ZN (n_3454), .A (n_3455));
NOR2_X1 i_2647 (.ZN (n_3453), .A1 (n_3462), .A2 (n_3454));
OAI21_X1 i_2646 (.ZN (n_3452), .A (n_3456), .B1 (n_3462), .B2 (n_3454));
XNOR2_X1 i_2645 (.ZN (n_3451), .A (n_3457), .B (n_3452));
NOR2_X1 i_2644 (.ZN (n_3450), .A1 (n_3486), .A2 (n_3451));
OAI21_X1 i_2643 (.ZN (n_3449), .A (n_3482), .B1 (n_3485), .B2 (n_3484));
NAND2_X1 i_2642 (.ZN (n_1750), .A1 (n_3483), .A2 (n_3449));
NOR2_X1 i_2641 (.ZN (n_3448), .A1 (n_3461), .A2 (n_3460));
XOR2_X1 i_2640 (.Z (n_1740), .A (n_3458), .B (n_3448));
NAND2_X1 i_2639 (.ZN (n_3447), .A1 (n_3481), .A2 (n_3471));
OAI21_X1 i_2638 (.ZN (n_1742), .A (n_3447), .B1 (n_3470), .B2 (n_3464));
FA_X1 i_2637 (.CO (n_1739), .S (n_3446), .A (n_1750), .B (n_1740), .CI (n_1742));
INV_X1 i_2636 (.ZN (n_3445), .A (inputB[31]));
INV_X2 i_2635 (.ZN (n_3444), .A (inputB[30]));
INV_X2 i_2634 (.ZN (n_3443), .A (inputB[29]));
INV_X2 i_2633 (.ZN (n_3442), .A (inputB[28]));
INV_X2 i_2632 (.ZN (n_3441), .A (inputB[27]));
INV_X2 i_2631 (.ZN (n_3440), .A (inputB[26]));
INV_X2 i_2630 (.ZN (n_3439), .A (inputB[25]));
INV_X2 i_2629 (.ZN (n_3438), .A (inputB[24]));
INV_X2 i_2628 (.ZN (n_3437), .A (inputB[23]));
INV_X2 i_2627 (.ZN (n_3436), .A (inputB[22]));
INV_X2 i_2626 (.ZN (n_3435), .A (inputB[21]));
INV_X2 i_2625 (.ZN (n_3434), .A (inputB[20]));
INV_X2 i_2624 (.ZN (n_3433), .A (inputB[19]));
INV_X2 i_2623 (.ZN (n_3432), .A (inputB[18]));
INV_X2 i_2622 (.ZN (n_3431), .A (inputB[17]));
INV_X2 i_2621 (.ZN (n_3430), .A (inputB[16]));
INV_X2 i_2620 (.ZN (n_3429), .A (inputB[15]));
INV_X2 i_2619 (.ZN (n_3428), .A (inputB[14]));
INV_X2 i_2618 (.ZN (n_3427), .A (inputB[13]));
INV_X2 i_2617 (.ZN (n_3426), .A (inputB[12]));
INV_X2 i_2616 (.ZN (n_3422), .A (inputB[11]));
INV_X2 i_2615 (.ZN (n_3421), .A (inputB[10]));
INV_X2 i_2614 (.ZN (n_3420), .A (inputB[9]));
INV_X2 i_2613 (.ZN (n_3419), .A (inputB[8]));
INV_X2 i_2612 (.ZN (n_3418), .A (inputB[7]));
INV_X2 i_2611 (.ZN (n_3417), .A (inputB[6]));
INV_X2 i_2610 (.ZN (n_3416), .A (inputB[5]));
INV_X2 i_2609 (.ZN (n_3415), .A (inputB[4]));
INV_X2 i_2608 (.ZN (n_3414), .A (inputB[3]));
INV_X4 i_2607 (.ZN (n_3413), .A (inputB[2]));
INV_X4 i_2606 (.ZN (n_3412), .A (inputB[1]));
INV_X2 i_2605 (.ZN (n_3411), .A (inputB[0]));
INV_X1 i_2604 (.ZN (n_3410), .A (inputA[31]));
INV_X1 i_2603 (.ZN (n_3406), .A (inputA[30]));
INV_X2 i_2602 (.ZN (n_3405), .A (inputA[29]));
INV_X2 i_2601 (.ZN (n_3404), .A (inputA[28]));
INV_X2 i_2600 (.ZN (n_2172), .A (inputA[27]));
INV_X2 i_2599 (.ZN (n_2171), .A (inputA[26]));
INV_X2 i_2598 (.ZN (n_2170), .A (inputA[25]));
INV_X2 i_2597 (.ZN (n_2169), .A (inputA[24]));
INV_X2 i_2596 (.ZN (n_2166), .A (inputA[23]));
INV_X2 i_2595 (.ZN (n_2164), .A (inputA[22]));
INV_X2 i_2594 (.ZN (n_2163), .A (inputA[21]));
INV_X2 i_2593 (.ZN (n_2162), .A (inputA[20]));
INV_X2 i_2592 (.ZN (n_2158), .A (inputA[19]));
INV_X2 i_2591 (.ZN (n_2156), .A (inputA[18]));
INV_X2 i_2590 (.ZN (n_2155), .A (inputA[17]));
INV_X2 i_2589 (.ZN (n_2154), .A (inputA[16]));
INV_X2 i_2588 (.ZN (n_2152), .A (inputA[15]));
INV_X2 i_2587 (.ZN (n_2151), .A (inputA[14]));
INV_X2 i_2586 (.ZN (n_2150), .A (inputA[13]));
INV_X2 i_2585 (.ZN (n_2149), .A (inputA[12]));
INV_X2 i_2584 (.ZN (n_2148), .A (inputA[11]));
INV_X2 i_2583 (.ZN (n_2146), .A (inputA[10]));
INV_X2 i_2582 (.ZN (n_2144), .A (inputA[9]));
INV_X2 i_2581 (.ZN (n_2143), .A (inputA[8]));
INV_X2 i_2580 (.ZN (n_2142), .A (inputA[7]));
INV_X2 i_2579 (.ZN (n_2141), .A (inputA[6]));
INV_X2 i_2578 (.ZN (n_2138), .A (inputA[5]));
INV_X2 i_2577 (.ZN (n_2136), .A (inputA[4]));
INV_X2 i_2576 (.ZN (n_2135), .A (inputA[3]));
INV_X2 i_2575 (.ZN (n_2134), .A (inputA[2]));
INV_X2 i_2574 (.ZN (n_2133), .A (inputA[1]));
NOR2_X1 i_2573 (.ZN (n_2132), .A1 (n_3443), .A2 (n_2138));
NAND2_X1 i_2572 (.ZN (n_2129), .A1 (inputB[31]), .A2 (inputA[3]));
NOR2_X1 i_2571 (.ZN (n_2128), .A1 (n_3444), .A2 (n_2136));
NAND2_X1 i_2570 (.ZN (n_2127), .A1 (n_2129), .A2 (n_2128));
NOR2_X1 i_2569 (.ZN (n_2126), .A1 (n_3445), .A2 (n_2133));
NAND2_X1 i_2568 (.ZN (n_2125), .A1 (inputB[30]), .A2 (inputA[2]));
NAND2_X1 i_2567 (.ZN (n_1777), .A1 (n_2126), .A2 (n_2125));
NAND2_X1 i_2566 (.ZN (n_1776), .A1 (inputB[31]), .A2 (inputA[0]));
NOR2_X1 i_2565 (.ZN (n_1775), .A1 (n_3444), .A2 (n_2133));
NAND2_X1 i_2564 (.ZN (n_1773), .A1 (n_1776), .A2 (n_1775));
NOR2_X1 i_2563 (.ZN (n_1772), .A1 (n_3443), .A2 (n_2134));
NAND2_X1 i_2562 (.ZN (n_1770), .A1 (inputB[31]), .A2 (inputA[2]));
NOR2_X1 i_2561 (.ZN (n_1769), .A1 (n_3444), .A2 (n_2135));
NAND2_X1 i_2560 (.ZN (n_1768), .A1 (n_1770), .A2 (n_1769));
NOR2_X1 i_2559 (.ZN (n_1767), .A1 (n_3443), .A2 (n_2136));
OAI211_X1 i_2558 (.ZN (n_1766), .A (inputB[0]), .B (inputA[31]), .C1 (n_3412), .C2 (n_3406));
AOI211_X1 i_2557 (.ZN (n_1763), .A (n_3412), .B (n_3406), .C1 (inputB[0]), .C2 (inputA[31]));
NAND2_X1 i_2556 (.ZN (n_1762), .A1 (inputB[4]), .A2 (inputA[30]));
NOR2_X1 i_2555 (.ZN (n_2926), .A1 (n_3414), .A2 (n_3405));
NOR3_X1 i_2554 (.ZN (n_1761), .A1 (n_3414), .A2 (n_3405), .A3 (n_1762));
AOI22_X1 i_2553 (.ZN (n_1759), .A1 (inputB[4]), .A2 (inputA[29]), .B1 (inputB[3]), .B2 (inputA[30]));
NOR2_X1 i_2552 (.ZN (n_1757), .A1 (n_3413), .A2 (n_3410));
OAI21_X1 i_2551 (.ZN (n_1756), .A (n_2127), .B1 (n_2129), .B2 (n_2128));
XNOR2_X1 i_2550 (.ZN (n_2124), .A (n_2132), .B (n_1756));
NOR2_X1 i_2549 (.ZN (n_2289), .A1 (n_3439), .A2 (n_2141));
NOR2_X1 i_2548 (.ZN (n_2318), .A1 (n_3438), .A2 (n_2142));
NOR2_X1 i_2547 (.ZN (n_2348), .A1 (n_3437), .A2 (n_2143));
NOR2_X1 i_2546 (.ZN (n_2202), .A1 (n_3442), .A2 (n_2135));
NOR2_X1 i_2545 (.ZN (n_2231), .A1 (n_3441), .A2 (n_2136));
NOR2_X1 i_2544 (.ZN (n_2261), .A1 (n_3440), .A2 (n_2138));
OAI21_X1 i_2543 (.ZN (n_1755), .A (n_1772), .B1 (n_1776), .B2 (n_1775));
NAND2_X1 i_2542 (.ZN (n_2165), .A1 (n_1773), .A2 (n_1755));
NOR2_X1 i_2541 (.ZN (n_2550), .A1 (n_3430), .A2 (n_2152));
NOR2_X1 i_2540 (.ZN (n_2579), .A1 (n_3429), .A2 (n_2154));
NOR2_X1 i_2539 (.ZN (n_2609), .A1 (n_3428), .A2 (n_2155));
NOR2_X1 i_2538 (.ZN (n_2463), .A1 (n_3433), .A2 (n_2149));
NOR2_X1 i_2537 (.ZN (n_2492), .A1 (n_3432), .A2 (n_2150));
NOR2_X1 i_2536 (.ZN (n_2522), .A1 (n_3431), .A2 (n_2151));
NOR2_X1 i_2535 (.ZN (n_2376), .A1 (n_3436), .A2 (n_2144));
NOR2_X1 i_2534 (.ZN (n_2405), .A1 (n_3435), .A2 (n_2146));
NOR2_X1 i_2533 (.ZN (n_2435), .A1 (n_3434), .A2 (n_2148));
NOR2_X1 i_2532 (.ZN (n_2287), .A1 (n_3439), .A2 (n_2143));
NOR2_X1 i_2531 (.ZN (n_2316), .A1 (n_3438), .A2 (n_2144));
NOR2_X1 i_2530 (.ZN (n_2346), .A1 (n_3437), .A2 (n_2146));
NOR2_X1 i_2529 (.ZN (n_2200), .A1 (n_3442), .A2 (n_2138));
NOR2_X1 i_2528 (.ZN (n_2229), .A1 (n_3441), .A2 (n_2141));
NOR2_X1 i_2527 (.ZN (n_2259), .A1 (n_3440), .A2 (n_2142));
OAI21_X1 i_2526 (.ZN (n_1754), .A (n_1767), .B1 (n_1770), .B2 (n_1769));
NAND2_X1 i_2525 (.ZN (n_2137), .A1 (n_1768), .A2 (n_1754));
NOR2_X1 i_2524 (.ZN (n_2811), .A1 (n_3418), .A2 (n_2169));
NOR2_X1 i_2523 (.ZN (n_2840), .A1 (n_3417), .A2 (n_2170));
NOR2_X1 i_2522 (.ZN (n_2870), .A1 (n_3416), .A2 (n_2171));
NOR2_X1 i_2521 (.ZN (n_2724), .A1 (n_3421), .A2 (n_2163));
NOR2_X1 i_2520 (.ZN (n_2753), .A1 (n_3420), .A2 (n_2164));
NOR2_X1 i_2519 (.ZN (n_2783), .A1 (n_3419), .A2 (n_2166));
NOR2_X1 i_2518 (.ZN (n_2637), .A1 (n_3427), .A2 (n_2156));
NOR2_X1 i_2517 (.ZN (n_2666), .A1 (n_3426), .A2 (n_2158));
NOR2_X1 i_2516 (.ZN (n_2696), .A1 (n_3422), .A2 (n_2162));
NOR2_X1 i_2515 (.ZN (n_2524), .A1 (n_3431), .A2 (n_2149));
NOR2_X1 i_2514 (.ZN (n_2552), .A1 (n_3430), .A2 (n_2150));
NOR2_X1 i_2513 (.ZN (n_2581), .A1 (n_3429), .A2 (n_2151));
NOR2_X1 i_2512 (.ZN (n_2437), .A1 (n_3434), .A2 (n_2144));
NOR2_X1 i_2511 (.ZN (n_2465), .A1 (n_3433), .A2 (n_2146));
NOR2_X1 i_2510 (.ZN (n_2494), .A1 (n_3432), .A2 (n_2148));
NOR2_X1 i_2509 (.ZN (n_2350), .A1 (n_3437), .A2 (n_2141));
NOR2_X1 i_2508 (.ZN (n_2378), .A1 (n_3436), .A2 (n_2142));
NOR2_X1 i_2507 (.ZN (n_2407), .A1 (n_3435), .A2 (n_2143));
NOR2_X1 i_2506 (.ZN (n_2785), .A1 (n_3419), .A2 (n_2163));
NOR2_X1 i_2505 (.ZN (n_2813), .A1 (n_3418), .A2 (n_2164));
NOR2_X1 i_2504 (.ZN (n_2842), .A1 (n_3417), .A2 (n_2166));
NOR2_X1 i_2503 (.ZN (n_2698), .A1 (n_3422), .A2 (n_2156));
NOR2_X1 i_2502 (.ZN (n_2726), .A1 (n_3421), .A2 (n_2158));
NOR2_X1 i_2501 (.ZN (n_2755), .A1 (n_3420), .A2 (n_2162));
NOR2_X1 i_2499 (.ZN (n_2611), .A1 (n_3428), .A2 (n_2152));
NOR2_X1 i_2498 (.ZN (n_2639), .A1 (n_3427), .A2 (n_2154));
NOR2_X1 i_2497 (.ZN (n_2668), .A1 (n_3426), .A2 (n_2155));
NOR2_X1 i_2496 (.ZN (n_3014), .A1 (n_3411), .A2 (n_3406));
NOR2_X1 i_2495 (.ZN (n_2958), .A1 (n_3413), .A2 (n_2172));
NOR2_X1 i_2493 (.ZN (n_2987), .A1 (n_3412), .A2 (n_3404));
NOR2_X1 i_2492 (.ZN (n_3015), .A1 (n_3411), .A2 (n_3405));
NOR2_X1 i_2491 (.ZN (n_2872), .A1 (n_3416), .A2 (n_2169));
NOR2_X1 i_2490 (.ZN (n_2900), .A1 (n_3415), .A2 (n_2170));
NOR2_X1 i_2489 (.ZN (n_2929), .A1 (n_3414), .A2 (n_2171));
NOR2_X1 i_2488 (.ZN (n_2782), .A1 (n_3419), .A2 (n_2169));
NOR2_X1 i_2487 (.ZN (n_2810), .A1 (n_3418), .A2 (n_2170));
NOR2_X1 i_2486 (.ZN (n_2839), .A1 (n_3417), .A2 (n_2171));
NOR2_X1 i_2485 (.ZN (n_2695), .A1 (n_3422), .A2 (n_2163));
NOR2_X1 i_2484 (.ZN (n_2723), .A1 (n_3421), .A2 (n_2164));
NOR2_X1 i_2483 (.ZN (n_2752), .A1 (n_3420), .A2 (n_2166));
NOR2_X1 i_2481 (.ZN (n_2608), .A1 (n_3428), .A2 (n_2156));
NOR2_X1 i_2480 (.ZN (n_2636), .A1 (n_3427), .A2 (n_2158));
NOR2_X1 i_2479 (.ZN (n_2665), .A1 (n_3426), .A2 (n_2162));
NOR2_X1 i_2478 (.ZN (n_2928), .A1 (n_3414), .A2 (n_2172));
NOR2_X1 i_2477 (.ZN (n_2957), .A1 (n_3413), .A2 (n_3404));
NOR2_X1 i_2476 (.ZN (n_2986), .A1 (n_3412), .A2 (n_3405));
OAI21_X1 i_2475 (.ZN (n_1751), .A (n_1766), .B1 (n_984), .B2 (n_1763));
INV_X1 i_2474 (.ZN (n_2157), .A (n_1751));
NOR2_X1 i_2473 (.ZN (n_2898), .A1 (n_3415), .A2 (n_2172));
NOR2_X1 i_2472 (.ZN (n_2927), .A1 (n_3414), .A2 (n_3404));
NOR2_X1 i_2471 (.ZN (n_2956), .A1 (n_3413), .A2 (n_3405));
NOR2_X1 i_2470 (.ZN (n_1749), .A1 (n_3412), .A2 (n_3410));
NOR3_X1 i_2469 (.ZN (n_1748), .A1 (n_3413), .A2 (n_3406), .A3 (n_1749));
OAI21_X1 i_2468 (.ZN (n_1747), .A (n_1749), .B1 (n_3413), .B2 (n_3406));
INV_X1 i_2467 (.ZN (n_1746), .A (n_1747));
NOR2_X1 i_2466 (.ZN (n_1744), .A1 (n_1748), .A2 (n_1746));
XOR2_X1 i_2465 (.Z (n_2147), .A (n_887), .B (n_1744));
NOR2_X1 i_2464 (.ZN (n_2869), .A1 (n_3416), .A2 (n_2172));
NOR2_X1 i_2463 (.ZN (n_2897), .A1 (n_3415), .A2 (n_3404));
OAI21_X1 i_2462 (.ZN (n_1741), .A (n_1747), .B1 (n_887), .B2 (n_1748));
INV_X1 i_2461 (.ZN (n_2145), .A (n_1741));
NOR2_X1 i_2460 (.ZN (n_1738), .A1 (n_1761), .A2 (n_1759));
XNOR2_X1 i_2459 (.ZN (n_2130), .A (n_1757), .B (n_1738));
FA_X1 i_2458 (.CO (n_1077), .S (n_1076), .A (n_1066), .B (n_1021), .CI (n_1019));
FA_X1 i_2457 (.CO (n_1019), .S (n_1067), .A (n_955), .B (n_953), .CI (n_1006));
FA_X1 i_2456 (.CO (n_1057), .S (n_1006), .A (n_945), .B (n_2145), .CI (n_2130));
FA_X1 i_2455 (.CO (n_953), .S (n_1020), .A (n_2157), .B (n_2147), .CI (n_942));
FA_X1 i_2454 (.CO (n_1018), .S (n_942), .A (n_2869), .B (n_2897), .CI (n_2926));
FA_X1 i_2453 (.CO (n_887), .S (n_1007), .A (n_2898), .B (n_2927), .CI (n_2956));
FA_X1 i_2452 (.CO (n_984), .S (n_982), .A (n_2928), .B (n_2957), .CI (n_2986));
FA_X1 i_2451 (.CO (n_955), .S (n_962), .A (n_940), .B (n_938), .CI (n_936));
FA_X1 i_2450 (.CO (n_960), .S (n_936), .A (n_2608), .B (n_2636), .CI (n_2665));
FA_X1 i_2449 (.CO (n_954), .S (n_938), .A (n_2695), .B (n_2723), .CI (n_2752));
FA_X1 i_2447 (.CO (n_952), .S (n_940), .A (n_2782), .B (n_2810), .CI (n_2839));
FA_X1 i_2445 (.CO (n_1021), .S (n_943), .A (n_1004), .B (n_963), .CI (n_961));
FA_X1 i_2444 (.CO (n_961), .S (n_941), .A (n_895), .B (n_948), .CI (n_946));
FA_X1 i_2443 (.CO (n_895), .S (n_939), .A (n_837), .B (n_835), .CI (n_833));
FA_X1 i_2442 (.CO (n_833), .S (n_937), .A (n_3014), .B (n_775), .CI (n_773));
FA_X1 i_2441 (.CO (n_773), .S (n_900), .A (n_2872), .B (n_2900), .CI (n_2929));
FA_X1 i_2440 (.CO (n_775), .S (n_898), .A (n_2958), .B (n_2987), .CI (n_3015));
FA_X1 i_2439 (.CO (n_835), .S (n_894), .A (n_771), .B (n_769), .CI (n_767));
FA_X1 i_2437 (.CO (n_767), .S (n_886), .A (n_2611), .B (n_2639), .CI (n_2668));
FA_X1 i_2436 (.CO (n_769), .S (n_884), .A (n_2698), .B (n_2726), .CI (n_2755));
FA_X1 i_2435 (.CO (n_771), .S (n_870), .A (n_2785), .B (n_2813), .CI (n_2842));
FA_X1 i_2434 (.CO (n_837), .S (n_836), .A (n_765), .B (n_763), .CI (n_761));
FA_X1 i_2433 (.CO (n_761), .S (n_834), .A (n_2350), .B (n_2378), .CI (n_2407));
FA_X1 i_2432 (.CO (n_763), .S (n_832), .A (n_2437), .B (n_2465), .CI (n_2494));
FA_X1 i_2430 (.CO (n_765), .S (n_831), .A (n_2524), .B (n_2552), .CI (n_2581));
FA_X1 i_2429 (.CO (n_963), .S (n_830), .A (n_944), .B (n_901), .CI (n_899));
FA_X1 i_2428 (.CO (n_899), .S (n_774), .A (n_882), .B (n_880), .CI (n_878));
FA_X1 i_2427 (.CO (n_901), .S (n_772), .A (n_876), .B (n_874), .CI (n_872));
FA_X1 i_2426 (.CO (n_945), .S (n_944), .A (n_885), .B (n_883), .CI (n_881));
FA_X1 i_2425 (.CO (n_881), .S (n_880), .A (n_2637), .B (n_2666), .CI (n_2696));
FA_X1 i_2424 (.CO (n_883), .S (n_882), .A (n_2724), .B (n_2753), .CI (n_2783));
FA_X1 i_2423 (.CO (n_885), .S (n_770), .A (n_2811), .B (n_2840), .CI (n_2870));
FA_X1 i_2422 (.CO (n_768), .S (n_1066), .A (n_2124), .B (n_1005), .CI (n_1056));
FA_X1 i_2421 (.CO (n_766), .S (n_1056), .A (n_985), .B (n_983), .CI (n_2137));
FA_X1 i_2420 (.CO (n_983), .S (n_764), .A (n_2200), .B (n_2229), .CI (n_2259));
FA_X1 i_2419 (.CO (n_985), .S (n_762), .A (n_2287), .B (n_2316), .CI (n_2346));
FA_X1 i_2418 (.CO (n_1005), .S (n_1004), .A (n_1777), .B (n_949), .CI (n_947));
FA_X1 i_2416 (.CO (n_947), .S (n_946), .A (n_879), .B (n_877), .CI (n_875));
FA_X1 i_2415 (.CO (n_875), .S (n_874), .A (n_2376), .B (n_2405), .CI (n_2435));
FA_X1 i_2414 (.CO (n_877), .S (n_876), .A (n_2463), .B (n_2492), .CI (n_2522));
FA_X1 i_2413 (.CO (n_879), .S (n_878), .A (n_2550), .B (n_2579), .CI (n_2609));
FA_X1 i_2412 (.CO (n_949), .S (n_948), .A (n_873), .B (n_871), .CI (n_2165));
FA_X1 i_2411 (.CO (n_871), .S (n_760), .A (n_2202), .B (n_2231), .CI (n_2261));
FA_X1 i_2410 (.CO (n_873), .S (n_872), .A (n_2289), .B (n_2318), .CI (n_2348));
INV_X2 i_2409 (.ZN (n_3425), .A (inputA[0]));
INV_X1 i_2408 (.ZN (n_3424), .A (n_925));
INV_X1 i_2407 (.ZN (n_3423), .A (n_980));
OAI21_X1 i_2406 (.ZN (n_3409), .A (n_3456), .B1 (n_3453), .B2 (n_3457));
INV_X1 i_2405 (.ZN (n_3408), .A (n_3409));
NOR2_X1 i_2404 (.ZN (n_3407), .A1 (n_3454), .A2 (n_3408));
AND2_X1 i_2403 (.ZN (n_3403), .A1 (n_6), .A2 (n_10));
NAND2_X1 i_2402 (.ZN (n_3402), .A1 (n_2), .A2 (n_4));
NOR2_X1 i_2401 (.ZN (n_3401), .A1 (n_3411), .A2 (n_2134));
NOR2_X1 i_2399 (.ZN (n_3400), .A1 (n_0), .A2 (n_3401));
NOR2_X1 i_2398 (.ZN (n_3399), .A1 (n_3412), .A2 (n_3425));
NOR2_X1 i_2397 (.ZN (n_3398), .A1 (n_3411), .A2 (n_2133));
NOR2_X1 i_2396 (.ZN (result[0]), .A1 (n_3411), .A2 (n_3425));
NOR2_X1 i_2395 (.ZN (n_3397), .A1 (n_3412), .A2 (n_2133));
NAND2_X1 i_2394 (.ZN (n_3396), .A1 (result[0]), .A2 (n_3397));
NAND2_X1 i_2393 (.ZN (n_3395), .A1 (n_0), .A2 (n_3401));
AOI21_X1 i_2392 (.ZN (n_3394), .A (n_3400), .B1 (n_3396), .B2 (n_3395));
OAI21_X1 i_2391 (.ZN (n_3393), .A (n_3394), .B1 (n_2), .B2 (n_4));
NAND2_X1 i_2390 (.ZN (n_3392), .A1 (n_3402), .A2 (n_3393));
OAI22_X1 i_2389 (.ZN (n_3391), .A1 (n_6), .A2 (n_10), .B1 (n_3403), .B2 (n_3392));
NOR2_X1 i_2388 (.ZN (n_3390), .A1 (n_52), .A2 (n_54));
NOR2_X1 i_2387 (.ZN (n_3389), .A1 (n_26), .A2 (n_28));
NOR2_X1 i_2385 (.ZN (n_3388), .A1 (n_38), .A2 (n_40));
OR3_X1 i_2384 (.ZN (n_3387), .A1 (n_3390), .A2 (n_3388), .A3 (n_3389));
NOR2_X1 i_2383 (.ZN (n_3386), .A1 (n_16), .A2 (n_18));
NOR3_X1 i_2382 (.ZN (n_3385), .A1 (n_3387), .A2 (n_3386), .A3 (n_3391));
NAND2_X1 i_2381 (.ZN (n_3384), .A1 (n_16), .A2 (n_18));
NAND2_X1 i_2380 (.ZN (n_3383), .A1 (n_26), .A2 (n_28));
AOI21_X1 i_2379 (.ZN (n_3382), .A (n_3387), .B1 (n_3384), .B2 (n_3383));
AND2_X1 i_2378 (.ZN (n_3381), .A1 (n_52), .A2 (n_54));
NAND2_X1 i_2377 (.ZN (n_3380), .A1 (n_38), .A2 (n_40));
INV_X1 i_2376 (.ZN (n_3379), .A (n_3380));
NOR2_X1 i_2375 (.ZN (n_3378), .A1 (n_3390), .A2 (n_3380));
NOR4_X1 i_2374 (.ZN (n_3377), .A1 (n_3381), .A2 (n_3378), .A3 (n_3382), .A4 (n_3385));
NOR2_X1 i_2373 (.ZN (n_3376), .A1 (n_128), .A2 (n_130));
NOR2_X1 i_2372 (.ZN (n_3375), .A1 (n_86), .A2 (n_88));
NOR2_X1 i_2371 (.ZN (n_3374), .A1 (n_106), .A2 (n_108));
OR3_X1 i_2370 (.ZN (n_3373), .A1 (n_3376), .A2 (n_3374), .A3 (n_3375));
NOR2_X1 i_2369 (.ZN (n_3372), .A1 (n_68), .A2 (n_70));
NOR3_X1 i_2368 (.ZN (n_3371), .A1 (n_3373), .A2 (n_3372), .A3 (n_3377));
NAND2_X1 i_2367 (.ZN (n_3370), .A1 (n_68), .A2 (n_70));
NAND2_X1 i_2366 (.ZN (n_3369), .A1 (n_86), .A2 (n_88));
AOI21_X1 i_2365 (.ZN (n_3368), .A (n_3373), .B1 (n_3370), .B2 (n_3369));
AND2_X1 i_2364 (.ZN (n_3367), .A1 (n_128), .A2 (n_130));
NAND2_X1 i_2363 (.ZN (n_3366), .A1 (n_106), .A2 (n_108));
INV_X1 i_2362 (.ZN (n_3365), .A (n_3366));
NOR2_X1 i_2361 (.ZN (n_3364), .A1 (n_3376), .A2 (n_3366));
NOR4_X1 i_2360 (.ZN (n_3363), .A1 (n_3367), .A2 (n_3364), .A3 (n_3368), .A4 (n_3371));
NOR2_X1 i_2358 (.ZN (n_3362), .A1 (n_236), .A2 (n_238));
NOR2_X1 i_2357 (.ZN (n_3361), .A1 (n_178), .A2 (n_180));
NOR2_X1 i_2355 (.ZN (n_3360), .A1 (n_206), .A2 (n_208));
OR3_X1 i_2323 (.ZN (n_3359), .A1 (n_3362), .A2 (n_3360), .A3 (n_3361));
NOR2_X1 i_2322 (.ZN (n_3358), .A1 (n_152), .A2 (n_154));
NOR3_X1 i_2321 (.ZN (n_3357), .A1 (n_3359), .A2 (n_3358), .A3 (n_3363));
NAND2_X1 i_2320 (.ZN (n_3356), .A1 (n_152), .A2 (n_154));
NAND2_X1 i_2319 (.ZN (n_3355), .A1 (n_178), .A2 (n_180));
AOI21_X1 i_2318 (.ZN (n_3354), .A (n_3359), .B1 (n_3356), .B2 (n_3355));
AND2_X1 i_2317 (.ZN (n_3353), .A1 (n_236), .A2 (n_238));
NAND2_X1 i_2316 (.ZN (n_3352), .A1 (n_206), .A2 (n_208));
INV_X1 i_2315 (.ZN (n_3351), .A (n_3352));
NOR2_X1 i_2314 (.ZN (n_3350), .A1 (n_3362), .A2 (n_3352));
NOR4_X2 i_2313 (.ZN (n_3349), .A1 (n_3353), .A2 (n_3350), .A3 (n_3354), .A4 (n_3357));
NOR2_X1 i_2312 (.ZN (n_3348), .A1 (n_379), .A2 (n_418));
NOR2_X1 i_2311 (.ZN (n_3347), .A1 (n_505), .A2 (n_550));
INV_X1 i_2310 (.ZN (n_3346), .A (n_3347));
NOR2_X1 i_2309 (.ZN (n_3345), .A1 (n_419), .A2 (n_460));
INV_X1 i_2308 (.ZN (n_3344), .A (n_3345));
NOR2_X1 i_2307 (.ZN (n_3343), .A1 (n_461), .A2 (n_504));
INV_X1 i_2269 (.ZN (n_3342), .A (n_3343));
NAND3_X1 i_2268 (.ZN (n_3341), .A1 (n_3346), .A2 (n_3342), .A3 (n_3344));
OR2_X1 i_2267 (.ZN (n_3340), .A1 (n_3348), .A2 (n_3341));
NOR2_X1 i_2266 (.ZN (n_3339), .A1 (n_925), .A2 (n_980));
INV_X1 i_2265 (.ZN (n_3338), .A (n_3339));
NOR2_X1 i_2264 (.ZN (n_3337), .A1 (n_811), .A2 (n_868));
INV_X1 i_2263 (.ZN (n_3336), .A (n_3337));
NOR2_X1 i_2261 (.ZN (n_3335), .A1 (n_869), .A2 (n_924));
INV_X1 i_2260 (.ZN (n_3334), .A (n_3335));
NAND3_X1 i_2259 (.ZN (n_3333), .A1 (n_3338), .A2 (n_3334), .A3 (n_3336));
NOR2_X1 i_2257 (.ZN (n_3332), .A1 (n_755), .A2 (n_810));
OR2_X1 i_2256 (.ZN (n_3331), .A1 (n_3333), .A2 (n_3332));
NOR2_X1 i_2226 (.ZN (n_3330), .A1 (n_701), .A2 (n_754));
INV_X1 i_2216 (.ZN (n_3329), .A (n_3330));
NOR2_X1 i_2215 (.ZN (n_3328), .A1 (n_599), .A2 (n_648));
INV_X1 i_2214 (.ZN (n_3327), .A (n_3328));
NOR2_X1 i_2213 (.ZN (n_3326), .A1 (n_649), .A2 (n_700));
INV_X1 i_2212 (.ZN (n_3325), .A (n_3326));
NAND3_X1 i_2211 (.ZN (n_3324), .A1 (n_3329), .A2 (n_3325), .A3 (n_3327));
NOR2_X1 i_2210 (.ZN (n_3323), .A1 (n_596), .A2 (n_598));
OR2_X1 i_2209 (.ZN (n_3322), .A1 (n_3324), .A2 (n_3323));
OR2_X1 i_2208 (.ZN (n_3321), .A1 (n_3331), .A2 (n_3322));
OR2_X1 i_2207 (.ZN (n_3320), .A1 (n_3340), .A2 (n_3321));
NOR2_X1 i_2206 (.ZN (n_3319), .A1 (n_376), .A2 (n_378));
INV_X1 i_2205 (.ZN (n_3318), .A (n_3319));
NOR2_X1 i_2204 (.ZN (n_3317), .A1 (n_271), .A2 (n_304));
INV_X1 i_2203 (.ZN (n_3316), .A (n_3317));
NOR2_X1 i_2202 (.ZN (n_3315), .A1 (n_305), .A2 (n_340));
INV_X1 i_2201 (.ZN (n_3314), .A (n_3315));
NAND3_X1 i_2200 (.ZN (n_3313), .A1 (n_3318), .A2 (n_3314), .A3 (n_3316));
NOR2_X1 i_2199 (.ZN (n_3312), .A1 (n_268), .A2 (n_270));
OR2_X1 i_2198 (.ZN (n_3311), .A1 (n_3313), .A2 (n_3312));
NOR3_X1 i_2197 (.ZN (n_3310), .A1 (n_3320), .A2 (n_3311), .A3 (n_3349));
NAND2_X1 i_2196 (.ZN (n_3309), .A1 (n_268), .A2 (n_270));
NAND2_X1 i_2195 (.ZN (n_3308), .A1 (n_271), .A2 (n_304));
INV_X1 i_2500 (.ZN (n_3307), .A (n_3308));
AOI21_X1 i_2194 (.ZN (n_3306), .A (n_3313), .B1 (n_3309), .B2 (n_3308));
AND2_X1 i_2193 (.ZN (n_3305), .A1 (n_305), .A2 (n_340));
AOI221_X1 i_2192 (.ZN (n_3304), .A (n_3306), .B1 (n_376), .B2 (n_378), .C1 (n_3318), .C2 (n_3305));
NAND2_X1 i_2191 (.ZN (n_3303), .A1 (n_596), .A2 (n_598));
NAND2_X1 i_2190 (.ZN (n_3302), .A1 (n_599), .A2 (n_648));
INV_X1 i_2494 (.ZN (n_3301), .A (n_3302));
AOI21_X1 i_2189 (.ZN (n_3300), .A (n_3324), .B1 (n_3303), .B2 (n_3302));
AND2_X1 i_2188 (.ZN (n_3299), .A1 (n_649), .A2 (n_700));
AOI221_X1 i_2187 (.ZN (n_3298), .A (n_3300), .B1 (n_701), .B2 (n_754), .C1 (n_3329), .C2 (n_3299));
NAND2_X1 i_2186 (.ZN (n_3297), .A1 (n_755), .A2 (n_810));
AND2_X1 i_2185 (.ZN (n_3296), .A1 (n_811), .A2 (n_868));
AOI21_X1 i_2184 (.ZN (n_3295), .A (n_3296), .B1 (n_755), .B2 (n_810));
NAND2_X1 i_2183 (.ZN (n_3294), .A1 (n_869), .A2 (n_924));
INV_X1 i_2182 (.ZN (n_3293), .A (n_3294));
OAI222_X1 i_2181 (.ZN (n_3292), .A1 (n_3333), .A2 (n_3295), .B1 (n_3339), .B2 (n_3294)
    , .C1 (n_3424), .C2 (n_3423));
NAND2_X1 i_2180 (.ZN (n_3291), .A1 (n_379), .A2 (n_418));
NAND2_X1 i_2179 (.ZN (n_3290), .A1 (n_419), .A2 (n_460));
INV_X1 i_2482 (.ZN (n_3289), .A (n_3290));
AOI21_X1 i_2178 (.ZN (n_3288), .A (n_3341), .B1 (n_3291), .B2 (n_3290));
AND2_X1 i_2177 (.ZN (n_3287), .A1 (n_461), .A2 (n_504));
AOI221_X1 i_2176 (.ZN (n_3286), .A (n_3288), .B1 (n_505), .B2 (n_550), .C1 (n_3346), .C2 (n_3287));
OAI222_X1 i_2175 (.ZN (n_3285), .A1 (n_3320), .A2 (n_3304), .B1 (n_3321), .B2 (n_3286)
    , .C1 (n_3331), .C2 (n_3298));
NOR3_X2 i_2174 (.ZN (n_3284), .A1 (n_3292), .A2 (n_3285), .A3 (n_3310));
NOR2_X1 i_2173 (.ZN (n_3283), .A1 (n_1185), .A2 (n_1230));
NOR2_X1 i_2172 (.ZN (n_3282), .A1 (n_1317), .A2 (n_1356));
INV_X1 i_2171 (.ZN (n_3281), .A (n_3282));
NOR2_X1 i_2170 (.ZN (n_3280), .A1 (n_1231), .A2 (n_1274));
INV_X1 i_2169 (.ZN (n_3279), .A (n_3280));
NOR2_X1 i_2168 (.ZN (n_3278), .A1 (n_1275), .A2 (n_1316));
INV_X1 i_2167 (.ZN (n_3277), .A (n_3278));
NAND3_X1 i_2166 (.ZN (n_3276), .A1 (n_3281), .A2 (n_3277), .A3 (n_3279));
OR2_X1 i_2165 (.ZN (n_3275), .A1 (n_3283), .A2 (n_3276));
NOR2_X1 i_2164 (.ZN (n_3274), .A1 (n_1581), .A2 (n_1604));
NOR2_X1 i_2163 (.ZN (n_3273), .A1 (n_1527), .A2 (n_1554));
NOR2_X1 i_2162 (.ZN (n_3272), .A1 (n_1555), .A2 (n_1580));
NOR2_X1 i_2161 (.ZN (n_3271), .A1 (n_3273), .A2 (n_3272));
NOR3_X1 i_2160 (.ZN (n_3270), .A1 (n_3274), .A2 (n_3272), .A3 (n_3273));
OAI21_X1 i_2159 (.ZN (n_3269), .A (n_3270), .B1 (n_1497), .B2 (n_1526));
NOR2_X1 i_2158 (.ZN (n_3268), .A1 (n_1465), .A2 (n_1496));
INV_X1 i_2157 (.ZN (n_3267), .A (n_3268));
NOR2_X1 i_2156 (.ZN (n_3266), .A1 (n_1395), .A2 (n_1430));
INV_X1 i_2155 (.ZN (n_3265), .A (n_3266));
NOR2_X1 i_2154 (.ZN (n_3264), .A1 (n_1431), .A2 (n_1464));
INV_X1 i_2153 (.ZN (n_3263), .A (n_3264));
NAND3_X1 i_2152 (.ZN (n_3262), .A1 (n_3267), .A2 (n_3263), .A3 (n_3265));
NOR2_X1 i_2151 (.ZN (n_3261), .A1 (n_1357), .A2 (n_1394));
OR2_X1 i_2150 (.ZN (n_3260), .A1 (n_3262), .A2 (n_3261));
OR2_X1 i_2149 (.ZN (n_3259), .A1 (n_3269), .A2 (n_3260));
OR2_X1 i_2148 (.ZN (n_3258), .A1 (n_3275), .A2 (n_3259));
NOR2_X1 i_2147 (.ZN (n_3257), .A1 (n_1137), .A2 (n_1184));
INV_X1 i_2146 (.ZN (n_3256), .A (n_3257));
NOR2_X1 i_2448 (.ZN (n_3255), .A1 (n_1035), .A2 (n_1086));
INV_X1 i_2145 (.ZN (n_3254), .A (n_3255));
NOR2_X1 i_2446 (.ZN (n_3253), .A1 (n_1087), .A2 (n_1136));
INV_X1 i_2144 (.ZN (n_3252), .A (n_3253));
NAND3_X1 i_2143 (.ZN (n_3251), .A1 (n_3256), .A2 (n_3252), .A3 (n_3254));
NOR2_X1 i_2142 (.ZN (n_3250), .A1 (n_981), .A2 (n_1034));
OR2_X1 i_2141 (.ZN (n_3249), .A1 (n_3251), .A2 (n_3250));
NOR3_X1 i_2140 (.ZN (n_3248), .A1 (n_3258), .A2 (n_3249), .A3 (n_3284));
NAND2_X1 i_2139 (.ZN (n_3247), .A1 (n_981), .A2 (n_1034));
NAND2_X1 i_2138 (.ZN (n_3246), .A1 (n_1035), .A2 (n_1086));
INV_X1 i_2438 (.ZN (n_3245), .A (n_3246));
AOI21_X1 i_2137 (.ZN (n_3244), .A (n_3251), .B1 (n_3247), .B2 (n_3246));
AND2_X1 i_2136 (.ZN (n_3243), .A1 (n_1087), .A2 (n_1136));
AOI221_X1 i_2135 (.ZN (n_3242), .A (n_3244), .B1 (n_1137), .B2 (n_1184), .C1 (n_3256), .C2 (n_3243));
NOR2_X1 i_2134 (.ZN (n_3241), .A1 (n_3258), .A2 (n_3242));
NAND2_X1 i_2133 (.ZN (n_3240), .A1 (n_1185), .A2 (n_1230));
NAND2_X1 i_2132 (.ZN (n_3239), .A1 (n_1231), .A2 (n_1274));
INV_X1 i_2431 (.ZN (n_3238), .A (n_3239));
AOI21_X1 i_2131 (.ZN (n_3237), .A (n_3276), .B1 (n_3240), .B2 (n_3239));
AND2_X1 i_2130 (.ZN (n_3236), .A1 (n_1275), .A2 (n_1316));
AOI221_X1 i_2129 (.ZN (n_3235), .A (n_3237), .B1 (n_1317), .B2 (n_1356), .C1 (n_3281), .C2 (n_3236));
NAND2_X1 i_2128 (.ZN (n_3234), .A1 (n_1497), .A2 (n_1526));
INV_X1 i_2127 (.ZN (n_3233), .A (n_3234));
AND2_X1 i_2126 (.ZN (n_3232), .A1 (n_1527), .A2 (n_1554));
OAI21_X1 i_2125 (.ZN (n_3231), .A (n_3270), .B1 (n_3233), .B2 (n_3232));
NAND2_X1 i_2124 (.ZN (n_3230), .A1 (n_1555), .A2 (n_1580));
INV_X1 i_2123 (.ZN (n_3229), .A (n_3230));
OAI21_X1 i_2122 (.ZN (n_3228), .A (n_3231), .B1 (n_3274), .B2 (n_3230));
AOI21_X1 i_2121 (.ZN (n_3227), .A (n_3228), .B1 (n_1581), .B2 (n_1604));
NAND2_X1 i_2120 (.ZN (n_3226), .A1 (n_1357), .A2 (n_1394));
NAND2_X1 i_2119 (.ZN (n_3225), .A1 (n_1395), .A2 (n_1430));
INV_X1 i_2417 (.ZN (n_3224), .A (n_3225));
AOI21_X1 i_2118 (.ZN (n_3223), .A (n_3262), .B1 (n_3226), .B2 (n_3225));
AND2_X1 i_2117 (.ZN (n_3222), .A1 (n_1431), .A2 (n_1464));
AOI221_X1 i_2116 (.ZN (n_3221), .A (n_3223), .B1 (n_1465), .B2 (n_1496), .C1 (n_3267), .C2 (n_3222));
OAI221_X1 i_2115 (.ZN (n_3220), .A (n_3227), .B1 (n_3269), .B2 (n_3221), .C1 (n_3259), .C2 (n_3235));
NOR3_X2 i_2114 (.ZN (n_3219), .A1 (n_3241), .A2 (n_3220), .A3 (n_3248));
NOR2_X1 i_2113 (.ZN (n_3218), .A1 (n_1665), .A2 (n_1680));
NOR2_X1 i_2112 (.ZN (n_3217), .A1 (n_1627), .A2 (n_1646));
NOR2_X1 i_2111 (.ZN (n_3216), .A1 (n_1647), .A2 (n_1664));
OR3_X1 i_2110 (.ZN (n_3215), .A1 (n_3218), .A2 (n_3216), .A3 (n_3217));
NOR2_X1 i_2109 (.ZN (n_3214), .A1 (n_1605), .A2 (n_1626));
NOR3_X1 i_2108 (.ZN (n_3213), .A1 (n_3215), .A2 (n_3214), .A3 (n_3219));
NAND2_X1 i_2107 (.ZN (n_3212), .A1 (n_1605), .A2 (n_1626));
NAND2_X1 i_2106 (.ZN (n_3211), .A1 (n_1627), .A2 (n_1646));
AOI21_X1 i_2105 (.ZN (n_3210), .A (n_3215), .B1 (n_3212), .B2 (n_3211));
AND2_X1 i_2104 (.ZN (n_3209), .A1 (n_1665), .A2 (n_1680));
NAND2_X1 i_2103 (.ZN (n_3208), .A1 (n_1647), .A2 (n_1664));
INV_X1 i_2400 (.ZN (n_3207), .A (n_3208));
NOR2_X1 i_2102 (.ZN (n_3206), .A1 (n_3218), .A2 (n_3208));
NOR4_X1 i_2101 (.ZN (n_3205), .A1 (n_3209), .A2 (n_3206), .A3 (n_3210), .A4 (n_3213));
NOR2_X1 i_2100 (.ZN (n_3204), .A1 (n_1717), .A2 (n_1724));
NOR2_X1 i_2099 (.ZN (n_3203), .A1 (n_1695), .A2 (n_1706));
NOR2_X1 i_2098 (.ZN (n_3202), .A1 (n_1707), .A2 (n_1716));
OR3_X1 i_2097 (.ZN (n_3201), .A1 (n_3204), .A2 (n_3202), .A3 (n_3203));
NOR2_X1 i_2096 (.ZN (n_3200), .A1 (n_1681), .A2 (n_1694));
NOR3_X1 i_2095 (.ZN (n_3199), .A1 (n_3201), .A2 (n_3200), .A3 (n_3205));
NAND2_X1 i_2094 (.ZN (n_3198), .A1 (n_1681), .A2 (n_1694));
NAND2_X1 i_2093 (.ZN (n_3197), .A1 (n_1695), .A2 (n_1706));
AOI21_X1 i_2092 (.ZN (n_3196), .A (n_3201), .B1 (n_3198), .B2 (n_3197));
AND2_X1 i_2091 (.ZN (n_3195), .A1 (n_1717), .A2 (n_1724));
NAND2_X1 i_2090 (.ZN (n_3194), .A1 (n_1707), .A2 (n_1716));
INV_X1 i_2386 (.ZN (n_3193), .A (n_3194));
NOR2_X1 i_2089 (.ZN (n_3192), .A1 (n_3204), .A2 (n_3194));
NOR4_X2 i_2088 (.ZN (n_3191), .A1 (n_3195), .A2 (n_3192), .A3 (n_3196), .A4 (n_3199));
NOR2_X1 i_2087 (.ZN (n_3190), .A1 (n_1737), .A2 (n_3446));
NOR2_X1 i_2086 (.ZN (n_3189), .A1 (n_1731), .A2 (n_1734));
NOR2_X1 i_2085 (.ZN (n_3188), .A1 (n_1735), .A2 (n_1736));
NOR3_X1 i_2084 (.ZN (n_3187), .A1 (n_3190), .A2 (n_3188), .A3 (n_3189));
INV_X1 i_2083 (.ZN (n_3186), .A (n_3187));
NOR2_X1 i_2082 (.ZN (n_3185), .A1 (n_1725), .A2 (n_1730));
NOR3_X1 i_2081 (.ZN (n_3184), .A1 (n_3186), .A2 (n_3185), .A3 (n_3191));
NAND2_X1 i_2080 (.ZN (n_3183), .A1 (n_1725), .A2 (n_1730));
INV_X1 i_2079 (.ZN (n_3182), .A (n_3183));
AND2_X1 i_2078 (.ZN (n_3181), .A1 (n_1731), .A2 (n_1734));
OAI21_X1 i_2077 (.ZN (n_3180), .A (n_3187), .B1 (n_3182), .B2 (n_3181));
INV_X1 i_2076 (.ZN (n_3179), .A (n_3180));
AND2_X1 i_2075 (.ZN (n_3178), .A1 (n_1737), .A2 (n_3446));
NAND2_X1 i_2074 (.ZN (n_3177), .A1 (n_1735), .A2 (n_1736));
NOR2_X1 i_2073 (.ZN (n_3176), .A1 (n_3190), .A2 (n_3177));
OR4_X1 i_2072 (.ZN (n_3175), .A1 (n_3178), .A2 (n_3176), .A3 (n_3179), .A4 (n_3184));
NOR2_X1 i_2071 (.ZN (n_3174), .A1 (n_3450), .A2 (n_3175));
AOI21_X1 i_2070 (.ZN (n_3173), .A (n_3174), .B1 (n_3486), .B2 (n_3451));
OAI22_X1 i_2069 (.ZN (result[63]), .A1 (n_3455), .A2 (n_3409), .B1 (n_3407), .B2 (n_3173));
AOI21_X1 i_2068 (.ZN (n_3172), .A (n_3407), .B1 (n_3454), .B2 (n_3408));
XOR2_X1 i_2067 (.Z (result[62]), .A (n_3173), .B (n_3172));
AOI21_X1 i_2066 (.ZN (n_3171), .A (n_3450), .B1 (n_3486), .B2 (n_3451));
XOR2_X1 i_2065 (.Z (result[61]), .A (n_3175), .B (n_3171));
NOR2_X1 i_2064 (.ZN (n_3170), .A1 (n_3190), .A2 (n_3178));
OR2_X1 i_2359 (.ZN (n_3169), .A1 (n_3185), .A2 (n_3182));
AOI21_X1 i_2063 (.ZN (n_3168), .A (n_3185), .B1 (n_3191), .B2 (n_3183));
NOR2_X1 i_2062 (.ZN (n_3167), .A1 (n_3189), .A2 (n_3181));
NAND2_X1 i_2356 (.ZN (n_3166), .A1 (n_3177), .A2 (n_3167));
OAI21_X1 i_2061 (.ZN (n_3165), .A (n_3177), .B1 (n_3189), .B2 (n_3188));
OAI21_X1 i_2354 (.ZN (n_3164), .A (n_3165), .B1 (n_3168), .B2 (n_3166));
XNOR2_X1 i_2353 (.ZN (result[60]), .A (n_3170), .B (n_3164));
AOI21_X1 i_2352 (.ZN (n_3163), .A (n_3188), .B1 (n_1735), .B2 (n_1736));
OAI22_X1 i_2351 (.ZN (n_3162), .A1 (n_1731), .A2 (n_1734), .B1 (n_3181), .B2 (n_3168));
XNOR2_X1 i_2350 (.ZN (result[59]), .A (n_3163), .B (n_3162));
XOR2_X1 i_2349 (.Z (result[58]), .A (n_3168), .B (n_3167));
XOR2_X1 i_2348 (.Z (result[57]), .A (n_3191), .B (n_3169));
NOR2_X1 i_2347 (.ZN (n_3161), .A1 (n_3204), .A2 (n_3195));
OAI21_X1 i_2346 (.ZN (n_3160), .A (n_3198), .B1 (n_1681), .B2 (n_1694));
AOI21_X1 i_2345 (.ZN (n_3159), .A (n_3200), .B1 (n_3205), .B2 (n_3198));
INV_X1 i_2344 (.ZN (n_3158), .A (n_3159));
AOI21_X1 i_2343 (.ZN (n_3157), .A (n_3203), .B1 (n_3197), .B2 (n_3158));
AOI21_X1 i_2342 (.ZN (n_3156), .A (n_3203), .B1 (n_1695), .B2 (n_1706));
OAI22_X1 i_2341 (.ZN (n_3155), .A1 (n_1707), .A2 (n_1716), .B1 (n_3193), .B2 (n_3157));
XNOR2_X1 i_2340 (.ZN (result[56]), .A (n_3161), .B (n_3155));
NOR2_X1 i_2339 (.ZN (n_3154), .A1 (n_3202), .A2 (n_3193));
XOR2_X1 i_2338 (.Z (result[55]), .A (n_3157), .B (n_3154));
XOR2_X1 i_2337 (.Z (result[54]), .A (n_3159), .B (n_3156));
XOR2_X1 i_2336 (.Z (result[53]), .A (n_3205), .B (n_3160));
NOR2_X1 i_2335 (.ZN (n_3153), .A1 (n_3218), .A2 (n_3209));
OAI21_X1 i_2334 (.ZN (n_3152), .A (n_3212), .B1 (n_1605), .B2 (n_1626));
AOI21_X1 i_2333 (.ZN (n_3151), .A (n_3214), .B1 (n_3219), .B2 (n_3212));
INV_X1 i_2332 (.ZN (n_3150), .A (n_3151));
AOI21_X1 i_2331 (.ZN (n_3149), .A (n_3217), .B1 (n_3211), .B2 (n_3150));
AOI21_X1 i_2330 (.ZN (n_3148), .A (n_3217), .B1 (n_1627), .B2 (n_1646));
OAI22_X1 i_2329 (.ZN (n_3147), .A1 (n_1647), .A2 (n_1664), .B1 (n_3207), .B2 (n_3149));
XNOR2_X1 i_2328 (.ZN (result[52]), .A (n_3153), .B (n_3147));
NOR2_X1 i_2327 (.ZN (n_3146), .A1 (n_3216), .A2 (n_3207));
XOR2_X1 i_2326 (.Z (result[51]), .A (n_3149), .B (n_3146));
XOR2_X1 i_2325 (.Z (result[50]), .A (n_3151), .B (n_3148));
XOR2_X1 i_2324 (.Z (result[49]), .A (n_3219), .B (n_3152));
AOI21_X1 i_2060 (.ZN (n_3145), .A (n_3274), .B1 (n_1581), .B2 (n_1604));
OAI21_X1 i_2059 (.ZN (n_3144), .A (n_3242), .B1 (n_3284), .B2 (n_3249));
INV_X1 i_2058 (.ZN (n_3143), .A (n_3144));
OAI21_X1 i_2057 (.ZN (n_3142), .A (n_3235), .B1 (n_3275), .B2 (n_3143));
INV_X1 i_2056 (.ZN (n_3141), .A (n_3142));
OAI21_X1 i_2055 (.ZN (n_3140), .A (n_3221), .B1 (n_3260), .B2 (n_3141));
OAI21_X1 i_2054 (.ZN (n_3139), .A (n_3234), .B1 (n_1497), .B2 (n_1526));
OAI22_X1 i_2053 (.ZN (n_3138), .A1 (n_1497), .A2 (n_1526), .B1 (n_3233), .B2 (n_3140));
INV_X1 i_2052 (.ZN (n_3137), .A (n_3138));
NOR2_X1 i_2051 (.ZN (n_3136), .A1 (n_3273), .A2 (n_3232));
NAND3_X1 i_2050 (.ZN (n_3135), .A1 (n_3230), .A2 (n_3136), .A3 (n_3138));
OAI21_X1 i_2049 (.ZN (n_3134), .A (n_3135), .B1 (n_3271), .B2 (n_3229));
XNOR2_X1 i_2048 (.ZN (result[48]), .A (n_3145), .B (n_3134));
NOR2_X1 i_2047 (.ZN (n_3133), .A1 (n_3272), .A2 (n_3229));
OAI22_X1 i_2046 (.ZN (n_3132), .A1 (n_1527), .A2 (n_1554), .B1 (n_3232), .B2 (n_3137));
XNOR2_X1 i_2045 (.ZN (result[47]), .A (n_3133), .B (n_3132));
XOR2_X1 i_2044 (.Z (result[46]), .A (n_3137), .B (n_3136));
XNOR2_X1 i_2306 (.ZN (result[45]), .A (n_3140), .B (n_3139));
AOI21_X1 i_2305 (.ZN (n_3131), .A (n_3268), .B1 (n_1465), .B2 (n_1496));
OAI21_X1 i_2304 (.ZN (n_3130), .A (n_3226), .B1 (n_1357), .B2 (n_1394));
AOI21_X1 i_2303 (.ZN (n_3129), .A (n_3261), .B1 (n_3226), .B2 (n_3141));
OAI21_X1 i_2302 (.ZN (n_3128), .A (n_3265), .B1 (n_3224), .B2 (n_3129));
INV_X1 i_2301 (.ZN (n_3127), .A (n_3128));
NOR2_X1 i_2300 (.ZN (n_3126), .A1 (n_3266), .A2 (n_3224));
OAI21_X1 i_2299 (.ZN (n_3125), .A (n_3263), .B1 (n_3222), .B2 (n_3127));
XNOR2_X1 i_2298 (.ZN (result[44]), .A (n_3131), .B (n_3125));
NOR2_X1 i_2297 (.ZN (n_3124), .A1 (n_3264), .A2 (n_3222));
XOR2_X1 i_2296 (.Z (result[43]), .A (n_3127), .B (n_3124));
XOR2_X1 i_2295 (.Z (result[42]), .A (n_3129), .B (n_3126));
XOR2_X1 i_2294 (.Z (result[41]), .A (n_3141), .B (n_3130));
AOI21_X1 i_2293 (.ZN (n_3123), .A (n_3282), .B1 (n_1317), .B2 (n_1356));
OAI21_X1 i_2292 (.ZN (n_3122), .A (n_3240), .B1 (n_1185), .B2 (n_1230));
AOI21_X1 i_2291 (.ZN (n_3121), .A (n_3283), .B1 (n_3240), .B2 (n_3143));
OAI21_X1 i_2290 (.ZN (n_3120), .A (n_3279), .B1 (n_3238), .B2 (n_3121));
INV_X1 i_2289 (.ZN (n_3119), .A (n_3120));
NOR2_X1 i_2288 (.ZN (n_3118), .A1 (n_3280), .A2 (n_3238));
OAI21_X1 i_2287 (.ZN (n_3117), .A (n_3277), .B1 (n_3236), .B2 (n_3119));
XNOR2_X1 i_2286 (.ZN (result[40]), .A (n_3123), .B (n_3117));
NOR2_X1 i_2285 (.ZN (n_3116), .A1 (n_3278), .A2 (n_3236));
XOR2_X1 i_2284 (.Z (result[39]), .A (n_3119), .B (n_3116));
XOR2_X1 i_2283 (.Z (result[38]), .A (n_3121), .B (n_3118));
XOR2_X1 i_2282 (.Z (result[37]), .A (n_3143), .B (n_3122));
AOI21_X1 i_2281 (.ZN (n_3115), .A (n_3257), .B1 (n_1137), .B2 (n_1184));
OAI21_X1 i_2280 (.ZN (n_3114), .A (n_3247), .B1 (n_981), .B2 (n_1034));
AOI21_X1 i_2279 (.ZN (n_3113), .A (n_3250), .B1 (n_3284), .B2 (n_3247));
OAI21_X1 i_2278 (.ZN (n_3112), .A (n_3254), .B1 (n_3245), .B2 (n_3113));
INV_X1 i_2277 (.ZN (n_3111), .A (n_3112));
NOR2_X1 i_2276 (.ZN (n_3110), .A1 (n_3255), .A2 (n_3245));
OAI21_X1 i_2275 (.ZN (n_3109), .A (n_3252), .B1 (n_3243), .B2 (n_3111));
XNOR2_X1 i_2274 (.ZN (result[36]), .A (n_3115), .B (n_3109));
NOR2_X1 i_2273 (.ZN (n_3108), .A1 (n_3253), .A2 (n_3243));
XOR2_X1 i_2272 (.Z (result[35]), .A (n_3111), .B (n_3108));
XOR2_X1 i_2271 (.Z (result[34]), .A (n_3113), .B (n_3110));
XOR2_X1 i_2270 (.Z (result[33]), .A (n_3284), .B (n_3114));
OAI21_X1 i_2043 (.ZN (n_3107), .A (n_3338), .B1 (n_3424), .B2 (n_3423));
OAI21_X1 i_2042 (.ZN (n_3106), .A (n_3304), .B1 (n_3349), .B2 (n_3311));
INV_X1 i_2041 (.ZN (n_3105), .A (n_3106));
OAI21_X1 i_2040 (.ZN (n_3104), .A (n_3286), .B1 (n_3340), .B2 (n_3105));
INV_X1 i_2039 (.ZN (n_3103), .A (n_3104));
OAI21_X1 i_2038 (.ZN (n_3102), .A (n_3298), .B1 (n_3322), .B2 (n_3103));
INV_X1 i_2037 (.ZN (n_3101), .A (n_3102));
OAI21_X1 i_2262 (.ZN (n_3100), .A (n_3297), .B1 (n_755), .B2 (n_810));
AOI21_X1 i_2036 (.ZN (n_3099), .A (n_3332), .B1 (n_3297), .B2 (n_3101));
OAI21_X1 i_2035 (.ZN (n_3098), .A (n_3336), .B1 (n_3296), .B2 (n_3099));
INV_X1 i_2034 (.ZN (n_3097), .A (n_3098));
NOR2_X1 i_2258 (.ZN (n_3096), .A1 (n_3337), .A2 (n_3296));
OAI21_X1 i_2033 (.ZN (n_3095), .A (n_3334), .B1 (n_3293), .B2 (n_3097));
XOR2_X1 i_2032 (.Z (result[32]), .A (n_3107), .B (n_3095));
NOR2_X1 i_2255 (.ZN (n_3094), .A1 (n_3335), .A2 (n_3293));
XOR2_X1 i_2254 (.Z (result[31]), .A (n_3097), .B (n_3094));
XOR2_X1 i_2253 (.Z (result[30]), .A (n_3099), .B (n_3096));
XOR2_X1 i_2252 (.Z (result[29]), .A (n_3101), .B (n_3100));
AOI21_X1 i_2251 (.ZN (n_3093), .A (n_3330), .B1 (n_701), .B2 (n_754));
OAI21_X1 i_2250 (.ZN (n_3092), .A (n_3303), .B1 (n_596), .B2 (n_598));
AOI21_X1 i_2249 (.ZN (n_3091), .A (n_3323), .B1 (n_3303), .B2 (n_3103));
OAI21_X1 i_2248 (.ZN (n_3090), .A (n_3327), .B1 (n_3301), .B2 (n_3091));
INV_X1 i_2247 (.ZN (n_3089), .A (n_3090));
NOR2_X1 i_2246 (.ZN (n_3088), .A1 (n_3328), .A2 (n_3301));
OAI21_X1 i_2245 (.ZN (n_3087), .A (n_3325), .B1 (n_3299), .B2 (n_3089));
XNOR2_X1 i_2244 (.ZN (result[28]), .A (n_3093), .B (n_3087));
NOR2_X1 i_2243 (.ZN (n_3086), .A1 (n_3326), .A2 (n_3299));
XOR2_X1 i_2242 (.Z (result[27]), .A (n_3089), .B (n_3086));
XOR2_X1 i_2241 (.Z (result[26]), .A (n_3091), .B (n_3088));
XOR2_X1 i_2240 (.Z (result[25]), .A (n_3103), .B (n_3092));
AOI21_X1 i_2239 (.ZN (n_3085), .A (n_3347), .B1 (n_505), .B2 (n_550));
OAI21_X1 i_2238 (.ZN (n_3084), .A (n_3291), .B1 (n_379), .B2 (n_418));
AOI21_X1 i_2237 (.ZN (n_3083), .A (n_3348), .B1 (n_3291), .B2 (n_3105));
OAI21_X1 i_2236 (.ZN (n_3082), .A (n_3344), .B1 (n_3289), .B2 (n_3083));
INV_X1 i_2235 (.ZN (n_3081), .A (n_3082));
NOR2_X1 i_2234 (.ZN (n_3080), .A1 (n_3345), .A2 (n_3289));
OAI21_X1 i_2233 (.ZN (n_3079), .A (n_3342), .B1 (n_3287), .B2 (n_3081));
XNOR2_X1 i_2232 (.ZN (result[24]), .A (n_3085), .B (n_3079));
NOR2_X1 i_2231 (.ZN (n_3078), .A1 (n_3343), .A2 (n_3287));
XOR2_X1 i_2230 (.Z (result[23]), .A (n_3081), .B (n_3078));
XOR2_X1 i_2229 (.Z (result[22]), .A (n_3083), .B (n_3080));
XOR2_X1 i_2228 (.Z (result[21]), .A (n_3105), .B (n_3084));
AOI21_X1 i_2227 (.ZN (n_3077), .A (n_3319), .B1 (n_376), .B2 (n_378));
OAI21_X1 i_2031 (.ZN (n_3076), .A (n_3309), .B1 (n_268), .B2 (n_270));
AOI21_X1 i_2225 (.ZN (n_3075), .A (n_3312), .B1 (n_3349), .B2 (n_3309));
OAI21_X1 i_2224 (.ZN (n_3074), .A (n_3316), .B1 (n_3307), .B2 (n_3075));
INV_X1 i_2223 (.ZN (n_3073), .A (n_3074));
NOR2_X1 i_2222 (.ZN (n_3072), .A1 (n_3317), .A2 (n_3307));
OAI21_X1 i_2221 (.ZN (n_3071), .A (n_3314), .B1 (n_3305), .B2 (n_3073));
XNOR2_X1 i_2220 (.ZN (result[20]), .A (n_3077), .B (n_3071));
NOR2_X1 i_2219 (.ZN (n_3070), .A1 (n_3315), .A2 (n_3305));
XOR2_X1 i_2218 (.Z (result[19]), .A (n_3073), .B (n_3070));
XOR2_X1 i_2217 (.Z (result[18]), .A (n_3075), .B (n_3072));
XOR2_X1 i_2030 (.Z (result[17]), .A (n_3349), .B (n_3076));
NOR2_X1 i_2029 (.ZN (n_3069), .A1 (n_3362), .A2 (n_3353));
OAI21_X1 i_2028 (.ZN (n_3068), .A (n_3356), .B1 (n_152), .B2 (n_154));
AOI21_X1 i_2027 (.ZN (n_3067), .A (n_3358), .B1 (n_3363), .B2 (n_3356));
INV_X1 i_2026 (.ZN (n_3066), .A (n_3067));
AOI21_X1 i_2025 (.ZN (n_3065), .A (n_3361), .B1 (n_3355), .B2 (n_3066));
AOI21_X1 i_2024 (.ZN (n_3064), .A (n_3361), .B1 (n_178), .B2 (n_180));
OAI22_X1 i_2023 (.ZN (n_3063), .A1 (n_206), .A2 (n_208), .B1 (n_3351), .B2 (n_3065));
XNOR2_X1 i_2022 (.ZN (result[16]), .A (n_3069), .B (n_3063));
NOR2_X1 i_2021 (.ZN (n_3062), .A1 (n_3360), .A2 (n_3351));
XOR2_X1 i_2020 (.Z (result[15]), .A (n_3065), .B (n_3062));
XOR2_X1 i_2019 (.Z (result[14]), .A (n_3067), .B (n_3064));
XOR2_X1 i_2018 (.Z (result[13]), .A (n_3363), .B (n_3068));
NOR2_X1 i_2017 (.ZN (n_3061), .A1 (n_3376), .A2 (n_3367));
OAI21_X1 i_2016 (.ZN (n_3060), .A (n_3370), .B1 (n_68), .B2 (n_70));
AOI21_X1 i_2015 (.ZN (n_3059), .A (n_3372), .B1 (n_3377), .B2 (n_3370));
INV_X1 i_2014 (.ZN (n_3058), .A (n_3059));
AOI21_X1 i_2013 (.ZN (n_3057), .A (n_3375), .B1 (n_3369), .B2 (n_3058));
AOI21_X1 i_2012 (.ZN (n_3056), .A (n_3375), .B1 (n_86), .B2 (n_88));
OAI22_X1 i_2011 (.ZN (n_3055), .A1 (n_106), .A2 (n_108), .B1 (n_3365), .B2 (n_3057));
XNOR2_X1 i_2010 (.ZN (result[12]), .A (n_3061), .B (n_3055));
NOR2_X1 i_2009 (.ZN (n_3054), .A1 (n_3374), .A2 (n_3365));
XOR2_X1 i_2008 (.Z (result[11]), .A (n_3057), .B (n_3054));
XOR2_X1 i_2007 (.Z (result[10]), .A (n_3059), .B (n_3056));
XOR2_X1 i_2006 (.Z (result[9]), .A (n_3377), .B (n_3060));
NOR2_X1 i_2005 (.ZN (n_3053), .A1 (n_3390), .A2 (n_3381));
OAI21_X1 i_2004 (.ZN (n_3052), .A (n_3384), .B1 (n_16), .B2 (n_18));
AOI21_X1 i_2003 (.ZN (n_3051), .A (n_3386), .B1 (n_3391), .B2 (n_3384));
INV_X1 i_2002 (.ZN (n_3050), .A (n_3051));
AOI21_X1 i_2001 (.ZN (n_3049), .A (n_3389), .B1 (n_3383), .B2 (n_3050));
AOI21_X1 i_2000 (.ZN (n_3048), .A (n_3389), .B1 (n_26), .B2 (n_28));
OAI22_X1 i_1999 (.ZN (n_3047), .A1 (n_38), .A2 (n_40), .B1 (n_3379), .B2 (n_3049));
XNOR2_X1 i_1998 (.ZN (result[8]), .A (n_3053), .B (n_3047));
NOR2_X1 i_1997 (.ZN (n_3046), .A1 (n_3388), .A2 (n_3379));
XOR2_X1 i_1996 (.Z (result[7]), .A (n_3049), .B (n_3046));
XOR2_X1 i_1995 (.Z (result[6]), .A (n_3051), .B (n_3048));
XOR2_X1 i_1994 (.Z (result[5]), .A (n_3391), .B (n_3052));
XOR2_X1 i_1993 (.Z (n_3045), .A (n_6), .B (n_10));
XOR2_X1 i_1992 (.Z (result[4]), .A (n_3392), .B (n_3045));
OAI21_X1 i_1991 (.ZN (n_3044), .A (n_3402), .B1 (n_2), .B2 (n_4));
XNOR2_X1 i_1990 (.ZN (result[3]), .A (n_3394), .B (n_3044));
OAI21_X1 i_1989 (.ZN (n_3043), .A (n_3395), .B1 (n_0), .B2 (n_3401));
XOR2_X1 i_1988 (.Z (result[2]), .A (n_3396), .B (n_3043));
OAI21_X1 i_1987 (.ZN (n_3042), .A (n_3396), .B1 (n_3399), .B2 (n_3398));
INV_X1 i_1986 (.ZN (result[1]), .A (n_3042));
NOR2_X1 i_1985 (.ZN (n_3041), .A1 (n_3411), .A2 (n_2135));
NOR2_X1 i_1984 (.ZN (n_3040), .A1 (n_3411), .A2 (n_2136));
NOR2_X1 i_1983 (.ZN (n_3039), .A1 (n_3411), .A2 (n_2138));
NOR2_X1 i_1982 (.ZN (n_3038), .A1 (n_3411), .A2 (n_2141));
NOR2_X1 i_1981 (.ZN (n_3037), .A1 (n_3411), .A2 (n_2142));
NOR2_X1 i_1980 (.ZN (n_3036), .A1 (n_3411), .A2 (n_2143));
NOR2_X1 i_1979 (.ZN (n_3035), .A1 (n_3411), .A2 (n_2144));
NOR2_X1 i_1978 (.ZN (n_3034), .A1 (n_3411), .A2 (n_2146));
NOR2_X1 i_1977 (.ZN (n_3033), .A1 (n_3411), .A2 (n_2148));
NOR2_X1 i_1976 (.ZN (n_3032), .A1 (n_3411), .A2 (n_2149));
NOR2_X1 i_1975 (.ZN (n_3031), .A1 (n_3411), .A2 (n_2150));
NOR2_X1 i_1974 (.ZN (n_3030), .A1 (n_3411), .A2 (n_2151));
NOR2_X1 i_1973 (.ZN (n_3029), .A1 (n_3411), .A2 (n_2152));
NOR2_X1 i_1972 (.ZN (n_3028), .A1 (n_3411), .A2 (n_2154));
NOR2_X1 i_1971 (.ZN (n_3027), .A1 (n_3411), .A2 (n_2155));
NOR2_X1 i_1970 (.ZN (n_3026), .A1 (n_3411), .A2 (n_2156));
NOR2_X1 i_1969 (.ZN (n_3025), .A1 (n_3411), .A2 (n_2158));
NOR2_X1 i_1968 (.ZN (n_3024), .A1 (n_3411), .A2 (n_2162));
NOR2_X1 i_1967 (.ZN (n_3023), .A1 (n_3411), .A2 (n_2163));
NOR2_X1 i_1966 (.ZN (n_3022), .A1 (n_3411), .A2 (n_2164));
NOR2_X1 i_1965 (.ZN (n_3021), .A1 (n_3411), .A2 (n_2166));
NOR2_X1 i_1964 (.ZN (n_3020), .A1 (n_3411), .A2 (n_2169));
NOR2_X1 i_1963 (.ZN (n_3019), .A1 (n_3411), .A2 (n_2170));
NOR2_X1 i_1962 (.ZN (n_3018), .A1 (n_3411), .A2 (n_2171));
NOR2_X1 i_1961 (.ZN (n_3017), .A1 (n_3411), .A2 (n_2172));
NOR2_X1 i_1960 (.ZN (n_3016), .A1 (n_3411), .A2 (n_3404));
NOR2_X1 i_1959 (.ZN (n_3013), .A1 (n_3412), .A2 (n_2134));
NOR2_X1 i_1958 (.ZN (n_3012), .A1 (n_3412), .A2 (n_2135));
NOR2_X1 i_1957 (.ZN (n_3011), .A1 (n_3412), .A2 (n_2136));
NOR2_X1 i_1956 (.ZN (n_3010), .A1 (n_3412), .A2 (n_2138));
NOR2_X1 i_1955 (.ZN (n_3009), .A1 (n_3412), .A2 (n_2141));
NOR2_X1 i_1954 (.ZN (n_3008), .A1 (n_3412), .A2 (n_2142));
NOR2_X1 i_1953 (.ZN (n_3007), .A1 (n_3412), .A2 (n_2143));
NOR2_X1 i_1952 (.ZN (n_3006), .A1 (n_3412), .A2 (n_2144));
NOR2_X1 i_1951 (.ZN (n_3005), .A1 (n_3412), .A2 (n_2146));
NOR2_X1 i_1950 (.ZN (n_3004), .A1 (n_3412), .A2 (n_2148));
NOR2_X1 i_1949 (.ZN (n_3003), .A1 (n_3412), .A2 (n_2149));
NOR2_X1 i_1948 (.ZN (n_3002), .A1 (n_3412), .A2 (n_2150));
NOR2_X1 i_1947 (.ZN (n_3001), .A1 (n_3412), .A2 (n_2151));
NOR2_X1 i_1946 (.ZN (n_3000), .A1 (n_3412), .A2 (n_2152));
NOR2_X1 i_1945 (.ZN (n_2999), .A1 (n_3412), .A2 (n_2154));
NOR2_X1 i_1944 (.ZN (n_2998), .A1 (n_3412), .A2 (n_2155));
NOR2_X1 i_1943 (.ZN (n_2997), .A1 (n_3412), .A2 (n_2156));
NOR2_X1 i_1942 (.ZN (n_2996), .A1 (n_3412), .A2 (n_2158));
NOR2_X1 i_1941 (.ZN (n_2995), .A1 (n_3412), .A2 (n_2162));
NOR2_X1 i_1940 (.ZN (n_2994), .A1 (n_3412), .A2 (n_2163));
NOR2_X1 i_1939 (.ZN (n_2993), .A1 (n_3412), .A2 (n_2164));
NOR2_X1 i_1938 (.ZN (n_2992), .A1 (n_3412), .A2 (n_2166));
NOR2_X1 i_1937 (.ZN (n_2991), .A1 (n_3412), .A2 (n_2169));
NOR2_X1 i_1936 (.ZN (n_2990), .A1 (n_3412), .A2 (n_2170));
NOR2_X1 i_1935 (.ZN (n_2989), .A1 (n_3412), .A2 (n_2171));
NOR2_X1 i_1934 (.ZN (n_2988), .A1 (n_3412), .A2 (n_2172));
NOR2_X1 i_1933 (.ZN (n_2985), .A1 (n_3413), .A2 (n_3425));
NOR2_X1 i_1932 (.ZN (n_2984), .A1 (n_3413), .A2 (n_2133));
NOR2_X1 i_1931 (.ZN (n_2983), .A1 (n_3413), .A2 (n_2134));
NOR2_X1 i_1930 (.ZN (n_2982), .A1 (n_3413), .A2 (n_2135));
NOR2_X1 i_1929 (.ZN (n_2981), .A1 (n_3413), .A2 (n_2136));
NOR2_X1 i_1928 (.ZN (n_2980), .A1 (n_3413), .A2 (n_2138));
NOR2_X1 i_1927 (.ZN (n_2979), .A1 (n_3413), .A2 (n_2141));
NOR2_X1 i_1926 (.ZN (n_2978), .A1 (n_3413), .A2 (n_2142));
NOR2_X1 i_1925 (.ZN (n_2977), .A1 (n_3413), .A2 (n_2143));
NOR2_X1 i_1924 (.ZN (n_2976), .A1 (n_3413), .A2 (n_2144));
NOR2_X1 i_1923 (.ZN (n_2975), .A1 (n_3413), .A2 (n_2146));
NOR2_X1 i_1922 (.ZN (n_2974), .A1 (n_3413), .A2 (n_2148));
NOR2_X1 i_1921 (.ZN (n_2973), .A1 (n_3413), .A2 (n_2149));
NOR2_X1 i_1920 (.ZN (n_2972), .A1 (n_3413), .A2 (n_2150));
NOR2_X1 i_1919 (.ZN (n_2971), .A1 (n_3413), .A2 (n_2151));
NOR2_X1 i_1918 (.ZN (n_2970), .A1 (n_3413), .A2 (n_2152));
NOR2_X1 i_1917 (.ZN (n_2969), .A1 (n_3413), .A2 (n_2154));
NOR2_X1 i_1916 (.ZN (n_2968), .A1 (n_3413), .A2 (n_2155));
NOR2_X1 i_1915 (.ZN (n_2967), .A1 (n_3413), .A2 (n_2156));
NOR2_X1 i_1914 (.ZN (n_2966), .A1 (n_3413), .A2 (n_2158));
NOR2_X1 i_1913 (.ZN (n_2965), .A1 (n_3413), .A2 (n_2162));
NOR2_X1 i_1912 (.ZN (n_2964), .A1 (n_3413), .A2 (n_2163));
NOR2_X1 i_1911 (.ZN (n_2963), .A1 (n_3413), .A2 (n_2164));
NOR2_X1 i_1910 (.ZN (n_2962), .A1 (n_3413), .A2 (n_2166));
NOR2_X1 i_1909 (.ZN (n_2961), .A1 (n_3413), .A2 (n_2169));
NOR2_X1 i_1908 (.ZN (n_2960), .A1 (n_3413), .A2 (n_2170));
NOR2_X1 i_1907 (.ZN (n_2959), .A1 (n_3413), .A2 (n_2171));
NOR2_X1 i_1906 (.ZN (n_2955), .A1 (n_3414), .A2 (n_3425));
NOR2_X1 i_1905 (.ZN (n_2954), .A1 (n_3414), .A2 (n_2133));
NOR2_X1 i_1904 (.ZN (n_2953), .A1 (n_3414), .A2 (n_2134));
NOR2_X1 i_1903 (.ZN (n_2952), .A1 (n_3414), .A2 (n_2135));
NOR2_X1 i_1902 (.ZN (n_2951), .A1 (n_3414), .A2 (n_2136));
NOR2_X1 i_1901 (.ZN (n_2950), .A1 (n_3414), .A2 (n_2138));
NOR2_X1 i_1900 (.ZN (n_2949), .A1 (n_3414), .A2 (n_2141));
NOR2_X1 i_1899 (.ZN (n_2948), .A1 (n_3414), .A2 (n_2142));
NOR2_X1 i_1898 (.ZN (n_2947), .A1 (n_3414), .A2 (n_2143));
NOR2_X1 i_1897 (.ZN (n_2946), .A1 (n_3414), .A2 (n_2144));
NOR2_X1 i_1896 (.ZN (n_2945), .A1 (n_3414), .A2 (n_2146));
NOR2_X1 i_1895 (.ZN (n_2944), .A1 (n_3414), .A2 (n_2148));
NOR2_X1 i_1894 (.ZN (n_2943), .A1 (n_3414), .A2 (n_2149));
NOR2_X1 i_1893 (.ZN (n_2942), .A1 (n_3414), .A2 (n_2150));
NOR2_X1 i_1892 (.ZN (n_2941), .A1 (n_3414), .A2 (n_2151));
NOR2_X1 i_1891 (.ZN (n_2940), .A1 (n_3414), .A2 (n_2152));
NOR2_X1 i_1890 (.ZN (n_2939), .A1 (n_3414), .A2 (n_2154));
NOR2_X1 i_1889 (.ZN (n_2938), .A1 (n_3414), .A2 (n_2155));
NOR2_X1 i_1888 (.ZN (n_2937), .A1 (n_3414), .A2 (n_2156));
NOR2_X1 i_1887 (.ZN (n_2936), .A1 (n_3414), .A2 (n_2158));
NOR2_X1 i_1886 (.ZN (n_2935), .A1 (n_3414), .A2 (n_2162));
NOR2_X1 i_1885 (.ZN (n_2934), .A1 (n_3414), .A2 (n_2163));
NOR2_X1 i_1884 (.ZN (n_2933), .A1 (n_3414), .A2 (n_2164));
NOR2_X1 i_1883 (.ZN (n_2932), .A1 (n_3414), .A2 (n_2166));
NOR2_X1 i_1882 (.ZN (n_2931), .A1 (n_3414), .A2 (n_2169));
NOR2_X1 i_1881 (.ZN (n_2930), .A1 (n_3414), .A2 (n_2170));
NOR2_X1 i_1880 (.ZN (n_2925), .A1 (n_3415), .A2 (n_3425));
NOR2_X1 i_1879 (.ZN (n_2924), .A1 (n_3415), .A2 (n_2133));
NOR2_X1 i_1878 (.ZN (n_2923), .A1 (n_3415), .A2 (n_2134));
NOR2_X1 i_1877 (.ZN (n_2922), .A1 (n_3415), .A2 (n_2135));
NOR2_X1 i_1876 (.ZN (n_2921), .A1 (n_3415), .A2 (n_2136));
NOR2_X1 i_1875 (.ZN (n_2920), .A1 (n_3415), .A2 (n_2138));
NOR2_X1 i_1874 (.ZN (n_2919), .A1 (n_3415), .A2 (n_2141));
NOR2_X1 i_1873 (.ZN (n_2918), .A1 (n_3415), .A2 (n_2142));
NOR2_X1 i_1872 (.ZN (n_2917), .A1 (n_3415), .A2 (n_2143));
NOR2_X1 i_1871 (.ZN (n_2916), .A1 (n_3415), .A2 (n_2144));
NOR2_X1 i_1870 (.ZN (n_2915), .A1 (n_3415), .A2 (n_2146));
NOR2_X1 i_1869 (.ZN (n_2914), .A1 (n_3415), .A2 (n_2148));
NOR2_X1 i_1868 (.ZN (n_2913), .A1 (n_3415), .A2 (n_2149));
NOR2_X1 i_1867 (.ZN (n_2912), .A1 (n_3415), .A2 (n_2150));
NOR2_X1 i_1866 (.ZN (n_2911), .A1 (n_3415), .A2 (n_2151));
NOR2_X1 i_1865 (.ZN (n_2910), .A1 (n_3415), .A2 (n_2152));
NOR2_X1 i_1864 (.ZN (n_2909), .A1 (n_3415), .A2 (n_2154));
NOR2_X1 i_1863 (.ZN (n_2908), .A1 (n_3415), .A2 (n_2155));
NOR2_X1 i_1862 (.ZN (n_2907), .A1 (n_3415), .A2 (n_2156));
NOR2_X1 i_1861 (.ZN (n_2906), .A1 (n_3415), .A2 (n_2158));
NOR2_X1 i_1860 (.ZN (n_2905), .A1 (n_3415), .A2 (n_2162));
NOR2_X1 i_1859 (.ZN (n_2904), .A1 (n_3415), .A2 (n_2163));
NOR2_X1 i_1858 (.ZN (n_2903), .A1 (n_3415), .A2 (n_2164));
NOR2_X1 i_1857 (.ZN (n_2902), .A1 (n_3415), .A2 (n_2166));
NOR2_X1 i_1856 (.ZN (n_2901), .A1 (n_3415), .A2 (n_2169));
NOR2_X1 i_1855 (.ZN (n_2899), .A1 (n_3415), .A2 (n_2171));
NOR2_X1 i_1854 (.ZN (n_2896), .A1 (n_3416), .A2 (n_3425));
NOR2_X1 i_1853 (.ZN (n_2895), .A1 (n_3416), .A2 (n_2133));
NOR2_X1 i_1852 (.ZN (n_2894), .A1 (n_3416), .A2 (n_2134));
NOR2_X1 i_1851 (.ZN (n_2893), .A1 (n_3416), .A2 (n_2135));
NOR2_X1 i_1850 (.ZN (n_2892), .A1 (n_3416), .A2 (n_2136));
NOR2_X1 i_1849 (.ZN (n_2891), .A1 (n_3416), .A2 (n_2138));
NOR2_X1 i_1848 (.ZN (n_2890), .A1 (n_3416), .A2 (n_2141));
NOR2_X1 i_1847 (.ZN (n_2889), .A1 (n_3416), .A2 (n_2142));
NOR2_X1 i_1846 (.ZN (n_2888), .A1 (n_3416), .A2 (n_2143));
NOR2_X1 i_1845 (.ZN (n_2887), .A1 (n_3416), .A2 (n_2144));
NOR2_X1 i_1844 (.ZN (n_2886), .A1 (n_3416), .A2 (n_2146));
NOR2_X1 i_1843 (.ZN (n_2885), .A1 (n_3416), .A2 (n_2148));
NOR2_X1 i_1842 (.ZN (n_2884), .A1 (n_3416), .A2 (n_2149));
NOR2_X1 i_1841 (.ZN (n_2883), .A1 (n_3416), .A2 (n_2150));
NOR2_X1 i_1840 (.ZN (n_2882), .A1 (n_3416), .A2 (n_2151));
NOR2_X1 i_1839 (.ZN (n_2881), .A1 (n_3416), .A2 (n_2152));
NOR2_X1 i_1838 (.ZN (n_2880), .A1 (n_3416), .A2 (n_2154));
NOR2_X1 i_1837 (.ZN (n_2879), .A1 (n_3416), .A2 (n_2155));
NOR2_X1 i_1836 (.ZN (n_2878), .A1 (n_3416), .A2 (n_2156));
NOR2_X1 i_1835 (.ZN (n_2877), .A1 (n_3416), .A2 (n_2158));
NOR2_X1 i_1834 (.ZN (n_2876), .A1 (n_3416), .A2 (n_2162));
NOR2_X1 i_1833 (.ZN (n_2875), .A1 (n_3416), .A2 (n_2163));
NOR2_X1 i_1832 (.ZN (n_2874), .A1 (n_3416), .A2 (n_2164));
NOR2_X1 i_1831 (.ZN (n_2873), .A1 (n_3416), .A2 (n_2166));
NOR2_X1 i_1830 (.ZN (n_2871), .A1 (n_3416), .A2 (n_2170));
NOR2_X1 i_1829 (.ZN (n_2868), .A1 (n_3416), .A2 (n_3404));
NOR2_X1 i_1828 (.ZN (n_2867), .A1 (n_3416), .A2 (n_3405));
NOR2_X1 i_1827 (.ZN (n_2866), .A1 (n_3416), .A2 (n_3406));
NOR2_X1 i_1826 (.ZN (n_2865), .A1 (n_3417), .A2 (n_3425));
NOR2_X1 i_1825 (.ZN (n_2864), .A1 (n_3417), .A2 (n_2133));
NOR2_X1 i_1824 (.ZN (n_2863), .A1 (n_3417), .A2 (n_2134));
NOR2_X1 i_1823 (.ZN (n_2862), .A1 (n_3417), .A2 (n_2135));
NOR2_X1 i_1822 (.ZN (n_2861), .A1 (n_3417), .A2 (n_2136));
NOR2_X1 i_1821 (.ZN (n_2860), .A1 (n_3417), .A2 (n_2138));
NOR2_X1 i_1820 (.ZN (n_2859), .A1 (n_3417), .A2 (n_2141));
NOR2_X1 i_1819 (.ZN (n_2858), .A1 (n_3417), .A2 (n_2142));
NOR2_X1 i_1818 (.ZN (n_2857), .A1 (n_3417), .A2 (n_2143));
NOR2_X1 i_1817 (.ZN (n_2856), .A1 (n_3417), .A2 (n_2144));
NOR2_X1 i_1816 (.ZN (n_2855), .A1 (n_3417), .A2 (n_2146));
NOR2_X1 i_1815 (.ZN (n_2854), .A1 (n_3417), .A2 (n_2148));
NOR2_X1 i_1814 (.ZN (n_2853), .A1 (n_3417), .A2 (n_2149));
NOR2_X1 i_1813 (.ZN (n_2852), .A1 (n_3417), .A2 (n_2150));
NOR2_X1 i_1812 (.ZN (n_2851), .A1 (n_3417), .A2 (n_2151));
NOR2_X1 i_1811 (.ZN (n_2850), .A1 (n_3417), .A2 (n_2152));
NOR2_X1 i_1810 (.ZN (n_2849), .A1 (n_3417), .A2 (n_2154));
NOR2_X1 i_1809 (.ZN (n_2848), .A1 (n_3417), .A2 (n_2155));
NOR2_X1 i_1808 (.ZN (n_2847), .A1 (n_3417), .A2 (n_2156));
NOR2_X1 i_1807 (.ZN (n_2846), .A1 (n_3417), .A2 (n_2158));
NOR2_X1 i_1806 (.ZN (n_2845), .A1 (n_3417), .A2 (n_2162));
NOR2_X1 i_1805 (.ZN (n_2844), .A1 (n_3417), .A2 (n_2163));
NOR2_X1 i_1804 (.ZN (n_2843), .A1 (n_3417), .A2 (n_2164));
NOR2_X1 i_1803 (.ZN (n_2841), .A1 (n_3417), .A2 (n_2169));
NOR2_X1 i_1802 (.ZN (n_2838), .A1 (n_3417), .A2 (n_2172));
NOR2_X1 i_1801 (.ZN (n_2837), .A1 (n_3417), .A2 (n_3404));
NOR2_X1 i_1800 (.ZN (n_2836), .A1 (n_3417), .A2 (n_3405));
NOR2_X1 i_1799 (.ZN (n_2835), .A1 (n_3418), .A2 (n_3425));
NOR2_X1 i_1798 (.ZN (n_2834), .A1 (n_3418), .A2 (n_2133));
NOR2_X1 i_1797 (.ZN (n_2833), .A1 (n_3418), .A2 (n_2134));
NOR2_X1 i_1796 (.ZN (n_2832), .A1 (n_3418), .A2 (n_2135));
NOR2_X1 i_1795 (.ZN (n_2831), .A1 (n_3418), .A2 (n_2136));
NOR2_X1 i_1794 (.ZN (n_2830), .A1 (n_3418), .A2 (n_2138));
NOR2_X1 i_1793 (.ZN (n_2829), .A1 (n_3418), .A2 (n_2141));
NOR2_X1 i_1792 (.ZN (n_2828), .A1 (n_3418), .A2 (n_2142));
NOR2_X1 i_1791 (.ZN (n_2827), .A1 (n_3418), .A2 (n_2143));
NOR2_X1 i_1790 (.ZN (n_2826), .A1 (n_3418), .A2 (n_2144));
NOR2_X1 i_1789 (.ZN (n_2825), .A1 (n_3418), .A2 (n_2146));
NOR2_X1 i_1788 (.ZN (n_2824), .A1 (n_3418), .A2 (n_2148));
NOR2_X1 i_1787 (.ZN (n_2823), .A1 (n_3418), .A2 (n_2149));
NOR2_X1 i_1786 (.ZN (n_2822), .A1 (n_3418), .A2 (n_2150));
NOR2_X1 i_1785 (.ZN (n_2821), .A1 (n_3418), .A2 (n_2151));
NOR2_X1 i_1784 (.ZN (n_2820), .A1 (n_3418), .A2 (n_2152));
NOR2_X1 i_1783 (.ZN (n_2819), .A1 (n_3418), .A2 (n_2154));
NOR2_X1 i_1782 (.ZN (n_2818), .A1 (n_3418), .A2 (n_2155));
NOR2_X1 i_1781 (.ZN (n_2817), .A1 (n_3418), .A2 (n_2156));
NOR2_X1 i_1780 (.ZN (n_2816), .A1 (n_3418), .A2 (n_2158));
NOR2_X1 i_1779 (.ZN (n_2815), .A1 (n_3418), .A2 (n_2162));
NOR2_X1 i_1778 (.ZN (n_2814), .A1 (n_3418), .A2 (n_2163));
NOR2_X1 i_1777 (.ZN (n_2812), .A1 (n_3418), .A2 (n_2166));
NOR2_X1 i_1776 (.ZN (n_2809), .A1 (n_3418), .A2 (n_2171));
NOR2_X1 i_1775 (.ZN (n_2808), .A1 (n_3418), .A2 (n_2172));
NOR2_X1 i_1774 (.ZN (n_2807), .A1 (n_3418), .A2 (n_3404));
NOR2_X1 i_1773 (.ZN (n_2806), .A1 (n_3419), .A2 (n_3425));
NOR2_X1 i_1772 (.ZN (n_2805), .A1 (n_3419), .A2 (n_2133));
NOR2_X1 i_1771 (.ZN (n_2804), .A1 (n_3419), .A2 (n_2134));
NOR2_X1 i_1770 (.ZN (n_2803), .A1 (n_3419), .A2 (n_2135));
NOR2_X1 i_1769 (.ZN (n_2802), .A1 (n_3419), .A2 (n_2136));
NOR2_X1 i_1768 (.ZN (n_2801), .A1 (n_3419), .A2 (n_2138));
NOR2_X1 i_1767 (.ZN (n_2800), .A1 (n_3419), .A2 (n_2141));
NOR2_X1 i_1766 (.ZN (n_2799), .A1 (n_3419), .A2 (n_2142));
NOR2_X1 i_1765 (.ZN (n_2798), .A1 (n_3419), .A2 (n_2143));
NOR2_X1 i_1764 (.ZN (n_2797), .A1 (n_3419), .A2 (n_2144));
NOR2_X1 i_1763 (.ZN (n_2796), .A1 (n_3419), .A2 (n_2146));
NOR2_X1 i_1762 (.ZN (n_2795), .A1 (n_3419), .A2 (n_2148));
NOR2_X1 i_1761 (.ZN (n_2794), .A1 (n_3419), .A2 (n_2149));
NOR2_X1 i_1760 (.ZN (n_2793), .A1 (n_3419), .A2 (n_2150));
NOR2_X1 i_1759 (.ZN (n_2792), .A1 (n_3419), .A2 (n_2151));
NOR2_X1 i_1758 (.ZN (n_2791), .A1 (n_3419), .A2 (n_2152));
NOR2_X1 i_1757 (.ZN (n_2790), .A1 (n_3419), .A2 (n_2154));
NOR2_X1 i_1756 (.ZN (n_2789), .A1 (n_3419), .A2 (n_2155));
NOR2_X1 i_1755 (.ZN (n_2788), .A1 (n_3419), .A2 (n_2156));
NOR2_X1 i_1754 (.ZN (n_2787), .A1 (n_3419), .A2 (n_2158));
NOR2_X1 i_1753 (.ZN (n_2786), .A1 (n_3419), .A2 (n_2162));
NOR2_X1 i_1752 (.ZN (n_2784), .A1 (n_3419), .A2 (n_2164));
NOR2_X1 i_1751 (.ZN (n_2781), .A1 (n_3419), .A2 (n_2170));
NOR2_X1 i_1750 (.ZN (n_2780), .A1 (n_3419), .A2 (n_2171));
NOR2_X1 i_1749 (.ZN (n_2779), .A1 (n_3419), .A2 (n_2172));
NOR2_X1 i_1748 (.ZN (n_2778), .A1 (n_3419), .A2 (n_3404));
NOR2_X1 i_1747 (.ZN (n_2777), .A1 (n_3419), .A2 (n_3405));
NOR2_X1 i_1746 (.ZN (n_2776), .A1 (n_3419), .A2 (n_3406));
NOR2_X1 i_1745 (.ZN (n_2775), .A1 (n_3420), .A2 (n_3425));
NOR2_X1 i_1744 (.ZN (n_2774), .A1 (n_3420), .A2 (n_2133));
NOR2_X1 i_1743 (.ZN (n_2773), .A1 (n_3420), .A2 (n_2134));
NOR2_X1 i_1742 (.ZN (n_2772), .A1 (n_3420), .A2 (n_2135));
NOR2_X1 i_1741 (.ZN (n_2771), .A1 (n_3420), .A2 (n_2136));
NOR2_X1 i_1740 (.ZN (n_2770), .A1 (n_3420), .A2 (n_2138));
NOR2_X1 i_1739 (.ZN (n_2769), .A1 (n_3420), .A2 (n_2141));
NOR2_X1 i_1738 (.ZN (n_2768), .A1 (n_3420), .A2 (n_2142));
NOR2_X1 i_1737 (.ZN (n_2767), .A1 (n_3420), .A2 (n_2143));
NOR2_X1 i_1736 (.ZN (n_2766), .A1 (n_3420), .A2 (n_2144));
NOR2_X1 i_1735 (.ZN (n_2765), .A1 (n_3420), .A2 (n_2146));
NOR2_X1 i_1734 (.ZN (n_2764), .A1 (n_3420), .A2 (n_2148));
NOR2_X1 i_1733 (.ZN (n_2763), .A1 (n_3420), .A2 (n_2149));
NOR2_X1 i_1732 (.ZN (n_2762), .A1 (n_3420), .A2 (n_2150));
NOR2_X1 i_1731 (.ZN (n_2761), .A1 (n_3420), .A2 (n_2151));
NOR2_X1 i_1730 (.ZN (n_2760), .A1 (n_3420), .A2 (n_2152));
NOR2_X1 i_1729 (.ZN (n_2759), .A1 (n_3420), .A2 (n_2154));
NOR2_X1 i_1728 (.ZN (n_2758), .A1 (n_3420), .A2 (n_2155));
NOR2_X1 i_1727 (.ZN (n_2757), .A1 (n_3420), .A2 (n_2156));
NOR2_X1 i_1726 (.ZN (n_2756), .A1 (n_3420), .A2 (n_2158));
NOR2_X1 i_1725 (.ZN (n_2754), .A1 (n_3420), .A2 (n_2163));
NOR2_X1 i_1724 (.ZN (n_2751), .A1 (n_3420), .A2 (n_2169));
NOR2_X1 i_1723 (.ZN (n_2750), .A1 (n_3420), .A2 (n_2170));
NOR2_X1 i_1722 (.ZN (n_2749), .A1 (n_3420), .A2 (n_2171));
NOR2_X1 i_1721 (.ZN (n_2748), .A1 (n_3420), .A2 (n_2172));
NOR2_X1 i_1720 (.ZN (n_2747), .A1 (n_3420), .A2 (n_3404));
NOR2_X1 i_1719 (.ZN (n_2746), .A1 (n_3420), .A2 (n_3405));
NOR2_X1 i_1718 (.ZN (n_2745), .A1 (n_3421), .A2 (n_3425));
NOR2_X1 i_1717 (.ZN (n_2744), .A1 (n_3421), .A2 (n_2133));
NOR2_X1 i_1716 (.ZN (n_2743), .A1 (n_3421), .A2 (n_2134));
NOR2_X1 i_1715 (.ZN (n_2742), .A1 (n_3421), .A2 (n_2135));
NOR2_X1 i_1714 (.ZN (n_2741), .A1 (n_3421), .A2 (n_2136));
NOR2_X1 i_1713 (.ZN (n_2740), .A1 (n_3421), .A2 (n_2138));
NOR2_X1 i_1712 (.ZN (n_2739), .A1 (n_3421), .A2 (n_2141));
NOR2_X1 i_1711 (.ZN (n_2738), .A1 (n_3421), .A2 (n_2142));
NOR2_X1 i_1710 (.ZN (n_2737), .A1 (n_3421), .A2 (n_2143));
NOR2_X1 i_1709 (.ZN (n_2736), .A1 (n_3421), .A2 (n_2144));
NOR2_X1 i_1708 (.ZN (n_2735), .A1 (n_3421), .A2 (n_2146));
NOR2_X1 i_1707 (.ZN (n_2734), .A1 (n_3421), .A2 (n_2148));
NOR2_X1 i_1706 (.ZN (n_2733), .A1 (n_3421), .A2 (n_2149));
NOR2_X1 i_1705 (.ZN (n_2732), .A1 (n_3421), .A2 (n_2150));
NOR2_X1 i_1704 (.ZN (n_2731), .A1 (n_3421), .A2 (n_2151));
NOR2_X1 i_1703 (.ZN (n_2730), .A1 (n_3421), .A2 (n_2152));
NOR2_X1 i_1702 (.ZN (n_2729), .A1 (n_3421), .A2 (n_2154));
NOR2_X1 i_1701 (.ZN (n_2728), .A1 (n_3421), .A2 (n_2155));
NOR2_X1 i_1700 (.ZN (n_2727), .A1 (n_3421), .A2 (n_2156));
NOR2_X1 i_1699 (.ZN (n_2725), .A1 (n_3421), .A2 (n_2162));
NOR2_X1 i_1698 (.ZN (n_2722), .A1 (n_3421), .A2 (n_2166));
NOR2_X1 i_1697 (.ZN (n_2721), .A1 (n_3421), .A2 (n_2169));
NOR2_X1 i_1696 (.ZN (n_2720), .A1 (n_3421), .A2 (n_2170));
NOR2_X1 i_1695 (.ZN (n_2719), .A1 (n_3421), .A2 (n_2171));
NOR2_X1 i_1694 (.ZN (n_2718), .A1 (n_3421), .A2 (n_2172));
NOR2_X1 i_1693 (.ZN (n_2717), .A1 (n_3421), .A2 (n_3404));
NOR2_X1 i_1692 (.ZN (n_2716), .A1 (n_3422), .A2 (n_3425));
NOR2_X1 i_1691 (.ZN (n_2715), .A1 (n_3422), .A2 (n_2133));
NOR2_X1 i_1690 (.ZN (n_2714), .A1 (n_3422), .A2 (n_2134));
NOR2_X1 i_1689 (.ZN (n_2713), .A1 (n_3422), .A2 (n_2135));
NOR2_X1 i_1688 (.ZN (n_2712), .A1 (n_3422), .A2 (n_2136));
NOR2_X1 i_1687 (.ZN (n_2711), .A1 (n_3422), .A2 (n_2138));
NOR2_X1 i_1686 (.ZN (n_2710), .A1 (n_3422), .A2 (n_2141));
NOR2_X1 i_1685 (.ZN (n_2709), .A1 (n_3422), .A2 (n_2142));
NOR2_X1 i_1684 (.ZN (n_2708), .A1 (n_3422), .A2 (n_2143));
NOR2_X1 i_1683 (.ZN (n_2707), .A1 (n_3422), .A2 (n_2144));
NOR2_X1 i_1682 (.ZN (n_2706), .A1 (n_3422), .A2 (n_2146));
NOR2_X1 i_1681 (.ZN (n_2705), .A1 (n_3422), .A2 (n_2148));
NOR2_X1 i_1680 (.ZN (n_2704), .A1 (n_3422), .A2 (n_2149));
NOR2_X1 i_1679 (.ZN (n_2703), .A1 (n_3422), .A2 (n_2150));
NOR2_X1 i_1678 (.ZN (n_2702), .A1 (n_3422), .A2 (n_2151));
NOR2_X1 i_1677 (.ZN (n_2701), .A1 (n_3422), .A2 (n_2152));
NOR2_X1 i_1676 (.ZN (n_2700), .A1 (n_3422), .A2 (n_2154));
NOR2_X1 i_1675 (.ZN (n_2699), .A1 (n_3422), .A2 (n_2155));
NOR2_X1 i_1674 (.ZN (n_2697), .A1 (n_3422), .A2 (n_2158));
NOR2_X1 i_1673 (.ZN (n_2694), .A1 (n_3422), .A2 (n_2164));
NOR2_X1 i_1672 (.ZN (n_2693), .A1 (n_3422), .A2 (n_2166));
NOR2_X1 i_1671 (.ZN (n_2692), .A1 (n_3422), .A2 (n_2169));
NOR2_X1 i_1670 (.ZN (n_2691), .A1 (n_3422), .A2 (n_2170));
NOR2_X1 i_1669 (.ZN (n_2690), .A1 (n_3422), .A2 (n_2171));
NOR2_X1 i_1668 (.ZN (n_2689), .A1 (n_3422), .A2 (n_2172));
NOR2_X1 i_1667 (.ZN (n_2688), .A1 (n_3422), .A2 (n_3404));
NOR2_X1 i_1666 (.ZN (n_2687), .A1 (n_3422), .A2 (n_3405));
NOR2_X1 i_1665 (.ZN (n_2686), .A1 (n_3422), .A2 (n_3406));
NOR2_X1 i_1664 (.ZN (n_2685), .A1 (n_3426), .A2 (n_3425));
NOR2_X1 i_1663 (.ZN (n_2684), .A1 (n_3426), .A2 (n_2133));
NOR2_X1 i_1662 (.ZN (n_2683), .A1 (n_3426), .A2 (n_2134));
NOR2_X1 i_1661 (.ZN (n_2682), .A1 (n_3426), .A2 (n_2135));
NOR2_X1 i_1660 (.ZN (n_2681), .A1 (n_3426), .A2 (n_2136));
NOR2_X1 i_1659 (.ZN (n_2680), .A1 (n_3426), .A2 (n_2138));
NOR2_X1 i_1658 (.ZN (n_2679), .A1 (n_3426), .A2 (n_2141));
NOR2_X1 i_1657 (.ZN (n_2678), .A1 (n_3426), .A2 (n_2142));
NOR2_X1 i_1656 (.ZN (n_2677), .A1 (n_3426), .A2 (n_2143));
NOR2_X1 i_1655 (.ZN (n_2676), .A1 (n_3426), .A2 (n_2144));
NOR2_X1 i_1654 (.ZN (n_2675), .A1 (n_3426), .A2 (n_2146));
NOR2_X1 i_1653 (.ZN (n_2674), .A1 (n_3426), .A2 (n_2148));
NOR2_X1 i_1652 (.ZN (n_2673), .A1 (n_3426), .A2 (n_2149));
NOR2_X1 i_1651 (.ZN (n_2672), .A1 (n_3426), .A2 (n_2150));
NOR2_X1 i_1650 (.ZN (n_2671), .A1 (n_3426), .A2 (n_2151));
NOR2_X1 i_1649 (.ZN (n_2670), .A1 (n_3426), .A2 (n_2152));
NOR2_X1 i_1648 (.ZN (n_2669), .A1 (n_3426), .A2 (n_2154));
NOR2_X1 i_1647 (.ZN (n_2667), .A1 (n_3426), .A2 (n_2156));
NOR2_X1 i_1646 (.ZN (n_2664), .A1 (n_3426), .A2 (n_2163));
NOR2_X1 i_1645 (.ZN (n_2663), .A1 (n_3426), .A2 (n_2164));
NOR2_X1 i_1644 (.ZN (n_2662), .A1 (n_3426), .A2 (n_2166));
NOR2_X1 i_1643 (.ZN (n_2661), .A1 (n_3426), .A2 (n_2169));
NOR2_X1 i_1642 (.ZN (n_2660), .A1 (n_3426), .A2 (n_2170));
NOR2_X1 i_1641 (.ZN (n_2659), .A1 (n_3426), .A2 (n_2171));
NOR2_X1 i_1640 (.ZN (n_2658), .A1 (n_3426), .A2 (n_2172));
NOR2_X1 i_1639 (.ZN (n_2657), .A1 (n_3426), .A2 (n_3404));
NOR2_X1 i_1638 (.ZN (n_2656), .A1 (n_3426), .A2 (n_3405));
NOR2_X1 i_1637 (.ZN (n_2655), .A1 (n_3427), .A2 (n_3425));
NOR2_X1 i_1636 (.ZN (n_2654), .A1 (n_3427), .A2 (n_2133));
NOR2_X1 i_1635 (.ZN (n_2653), .A1 (n_3427), .A2 (n_2134));
NOR2_X1 i_1634 (.ZN (n_2652), .A1 (n_3427), .A2 (n_2135));
NOR2_X1 i_1633 (.ZN (n_2651), .A1 (n_3427), .A2 (n_2136));
NOR2_X1 i_1632 (.ZN (n_2650), .A1 (n_3427), .A2 (n_2138));
NOR2_X1 i_1631 (.ZN (n_2649), .A1 (n_3427), .A2 (n_2141));
NOR2_X1 i_1630 (.ZN (n_2648), .A1 (n_3427), .A2 (n_2142));
NOR2_X1 i_1629 (.ZN (n_2647), .A1 (n_3427), .A2 (n_2143));
NOR2_X1 i_1628 (.ZN (n_2646), .A1 (n_3427), .A2 (n_2144));
NOR2_X1 i_1627 (.ZN (n_2645), .A1 (n_3427), .A2 (n_2146));
NOR2_X1 i_1626 (.ZN (n_2644), .A1 (n_3427), .A2 (n_2148));
NOR2_X1 i_1625 (.ZN (n_2643), .A1 (n_3427), .A2 (n_2149));
NOR2_X1 i_1624 (.ZN (n_2642), .A1 (n_3427), .A2 (n_2150));
NOR2_X1 i_1623 (.ZN (n_2641), .A1 (n_3427), .A2 (n_2151));
NOR2_X1 i_1622 (.ZN (n_2640), .A1 (n_3427), .A2 (n_2152));
NOR2_X1 i_1621 (.ZN (n_2638), .A1 (n_3427), .A2 (n_2155));
NOR2_X1 i_1620 (.ZN (n_2635), .A1 (n_3427), .A2 (n_2162));
NOR2_X1 i_1619 (.ZN (n_2634), .A1 (n_3427), .A2 (n_2163));
NOR2_X1 i_1618 (.ZN (n_2633), .A1 (n_3427), .A2 (n_2164));
NOR2_X1 i_1617 (.ZN (n_2632), .A1 (n_3427), .A2 (n_2166));
NOR2_X1 i_1616 (.ZN (n_2631), .A1 (n_3427), .A2 (n_2169));
NOR2_X1 i_1615 (.ZN (n_2630), .A1 (n_3427), .A2 (n_2170));
NOR2_X1 i_1614 (.ZN (n_2629), .A1 (n_3427), .A2 (n_2171));
NOR2_X1 i_1613 (.ZN (n_2628), .A1 (n_3427), .A2 (n_2172));
NOR2_X1 i_1612 (.ZN (n_2627), .A1 (n_3427), .A2 (n_3404));
NOR2_X1 i_1611 (.ZN (n_2626), .A1 (n_3428), .A2 (n_3425));
NOR2_X1 i_1610 (.ZN (n_2625), .A1 (n_3428), .A2 (n_2133));
NOR2_X1 i_1609 (.ZN (n_2624), .A1 (n_3428), .A2 (n_2134));
NOR2_X1 i_1608 (.ZN (n_2623), .A1 (n_3428), .A2 (n_2135));
NOR2_X1 i_1607 (.ZN (n_2622), .A1 (n_3428), .A2 (n_2136));
NOR2_X1 i_1606 (.ZN (n_2621), .A1 (n_3428), .A2 (n_2138));
NOR2_X1 i_1605 (.ZN (n_2620), .A1 (n_3428), .A2 (n_2141));
NOR2_X1 i_1604 (.ZN (n_2619), .A1 (n_3428), .A2 (n_2142));
NOR2_X1 i_1603 (.ZN (n_2618), .A1 (n_3428), .A2 (n_2143));
NOR2_X1 i_1602 (.ZN (n_2617), .A1 (n_3428), .A2 (n_2144));
NOR2_X1 i_1601 (.ZN (n_2616), .A1 (n_3428), .A2 (n_2146));
NOR2_X1 i_1600 (.ZN (n_2615), .A1 (n_3428), .A2 (n_2148));
NOR2_X1 i_1599 (.ZN (n_2614), .A1 (n_3428), .A2 (n_2149));
NOR2_X1 i_1598 (.ZN (n_2613), .A1 (n_3428), .A2 (n_2150));
NOR2_X1 i_1597 (.ZN (n_2612), .A1 (n_3428), .A2 (n_2151));
NOR2_X1 i_1596 (.ZN (n_2610), .A1 (n_3428), .A2 (n_2154));
NOR2_X1 i_1595 (.ZN (n_2607), .A1 (n_3428), .A2 (n_2158));
NOR2_X1 i_1594 (.ZN (n_2606), .A1 (n_3428), .A2 (n_2162));
NOR2_X1 i_1593 (.ZN (n_2605), .A1 (n_3428), .A2 (n_2163));
NOR2_X1 i_1592 (.ZN (n_2604), .A1 (n_3428), .A2 (n_2164));
NOR2_X1 i_1591 (.ZN (n_2603), .A1 (n_3428), .A2 (n_2166));
NOR2_X1 i_1590 (.ZN (n_2602), .A1 (n_3428), .A2 (n_2169));
NOR2_X1 i_1589 (.ZN (n_2601), .A1 (n_3428), .A2 (n_2170));
NOR2_X1 i_1588 (.ZN (n_2600), .A1 (n_3428), .A2 (n_2171));
NOR2_X1 i_1587 (.ZN (n_2599), .A1 (n_3428), .A2 (n_2172));
NOR2_X1 i_1586 (.ZN (n_2598), .A1 (n_3428), .A2 (n_3404));
NOR2_X1 i_1585 (.ZN (n_2597), .A1 (n_3428), .A2 (n_3405));
NOR2_X1 i_1584 (.ZN (n_2596), .A1 (n_3428), .A2 (n_3406));
NOR2_X1 i_1583 (.ZN (n_2595), .A1 (n_3429), .A2 (n_3425));
NOR2_X1 i_1582 (.ZN (n_2594), .A1 (n_3429), .A2 (n_2133));
NOR2_X1 i_1581 (.ZN (n_2593), .A1 (n_3429), .A2 (n_2134));
NOR2_X1 i_1580 (.ZN (n_2592), .A1 (n_3429), .A2 (n_2135));
NOR2_X1 i_1579 (.ZN (n_2591), .A1 (n_3429), .A2 (n_2136));
NOR2_X1 i_1578 (.ZN (n_2590), .A1 (n_3429), .A2 (n_2138));
NOR2_X1 i_1577 (.ZN (n_2589), .A1 (n_3429), .A2 (n_2141));
NOR2_X1 i_1576 (.ZN (n_2588), .A1 (n_3429), .A2 (n_2142));
NOR2_X1 i_1575 (.ZN (n_2587), .A1 (n_3429), .A2 (n_2143));
NOR2_X1 i_1574 (.ZN (n_2586), .A1 (n_3429), .A2 (n_2144));
NOR2_X1 i_1573 (.ZN (n_2585), .A1 (n_3429), .A2 (n_2146));
NOR2_X1 i_1572 (.ZN (n_2584), .A1 (n_3429), .A2 (n_2148));
NOR2_X1 i_1571 (.ZN (n_2583), .A1 (n_3429), .A2 (n_2149));
NOR2_X1 i_1570 (.ZN (n_2582), .A1 (n_3429), .A2 (n_2150));
NOR2_X1 i_1569 (.ZN (n_2580), .A1 (n_3429), .A2 (n_2152));
NOR2_X1 i_1568 (.ZN (n_2578), .A1 (n_3429), .A2 (n_2155));
NOR2_X1 i_1567 (.ZN (n_2577), .A1 (n_3429), .A2 (n_2156));
NOR2_X1 i_1566 (.ZN (n_2576), .A1 (n_3429), .A2 (n_2158));
NOR2_X1 i_1565 (.ZN (n_2575), .A1 (n_3429), .A2 (n_2162));
NOR2_X1 i_1564 (.ZN (n_2574), .A1 (n_3429), .A2 (n_2163));
NOR2_X1 i_1563 (.ZN (n_2573), .A1 (n_3429), .A2 (n_2164));
NOR2_X1 i_1562 (.ZN (n_2572), .A1 (n_3429), .A2 (n_2166));
NOR2_X1 i_1561 (.ZN (n_2571), .A1 (n_3429), .A2 (n_2169));
NOR2_X1 i_1560 (.ZN (n_2570), .A1 (n_3429), .A2 (n_2170));
NOR2_X1 i_1559 (.ZN (n_2569), .A1 (n_3429), .A2 (n_2171));
NOR2_X1 i_1558 (.ZN (n_2568), .A1 (n_3429), .A2 (n_2172));
NOR2_X1 i_1557 (.ZN (n_2567), .A1 (n_3429), .A2 (n_3404));
NOR2_X1 i_1556 (.ZN (n_2566), .A1 (n_3429), .A2 (n_3405));
NOR2_X1 i_1555 (.ZN (n_2565), .A1 (n_3430), .A2 (n_3425));
NOR2_X1 i_1554 (.ZN (n_2564), .A1 (n_3430), .A2 (n_2133));
NOR2_X1 i_1553 (.ZN (n_2563), .A1 (n_3430), .A2 (n_2134));
NOR2_X1 i_1552 (.ZN (n_2562), .A1 (n_3430), .A2 (n_2135));
NOR2_X1 i_1551 (.ZN (n_2561), .A1 (n_3430), .A2 (n_2136));
NOR2_X1 i_1550 (.ZN (n_2560), .A1 (n_3430), .A2 (n_2138));
NOR2_X1 i_1549 (.ZN (n_2559), .A1 (n_3430), .A2 (n_2141));
NOR2_X1 i_1548 (.ZN (n_2558), .A1 (n_3430), .A2 (n_2142));
NOR2_X1 i_1547 (.ZN (n_2557), .A1 (n_3430), .A2 (n_2143));
NOR2_X1 i_1546 (.ZN (n_2556), .A1 (n_3430), .A2 (n_2144));
NOR2_X1 i_1545 (.ZN (n_2555), .A1 (n_3430), .A2 (n_2146));
NOR2_X1 i_1544 (.ZN (n_2554), .A1 (n_3430), .A2 (n_2148));
NOR2_X1 i_1543 (.ZN (n_2553), .A1 (n_3430), .A2 (n_2149));
NOR2_X1 i_1542 (.ZN (n_2551), .A1 (n_3430), .A2 (n_2151));
NOR2_X1 i_1541 (.ZN (n_2549), .A1 (n_3430), .A2 (n_2154));
NOR2_X1 i_1540 (.ZN (n_2548), .A1 (n_3430), .A2 (n_2155));
NOR2_X1 i_1539 (.ZN (n_2547), .A1 (n_3430), .A2 (n_2156));
NOR2_X1 i_1538 (.ZN (n_2546), .A1 (n_3430), .A2 (n_2158));
NOR2_X1 i_1537 (.ZN (n_2545), .A1 (n_3430), .A2 (n_2162));
NOR2_X1 i_1536 (.ZN (n_2544), .A1 (n_3430), .A2 (n_2163));
NOR2_X1 i_1535 (.ZN (n_2543), .A1 (n_3430), .A2 (n_2164));
NOR2_X1 i_1534 (.ZN (n_2542), .A1 (n_3430), .A2 (n_2166));
NOR2_X1 i_1533 (.ZN (n_2541), .A1 (n_3430), .A2 (n_2169));
NOR2_X1 i_1532 (.ZN (n_2540), .A1 (n_3430), .A2 (n_2170));
NOR2_X1 i_1531 (.ZN (n_2539), .A1 (n_3430), .A2 (n_2171));
NOR2_X1 i_1530 (.ZN (n_2538), .A1 (n_3430), .A2 (n_2172));
NOR2_X1 i_1529 (.ZN (n_2537), .A1 (n_3430), .A2 (n_3404));
NOR2_X1 i_1528 (.ZN (n_2536), .A1 (n_3431), .A2 (n_3425));
NOR2_X1 i_1527 (.ZN (n_2535), .A1 (n_3431), .A2 (n_2133));
NOR2_X1 i_1526 (.ZN (n_2534), .A1 (n_3431), .A2 (n_2134));
NOR2_X1 i_1525 (.ZN (n_2533), .A1 (n_3431), .A2 (n_2135));
NOR2_X1 i_1524 (.ZN (n_2532), .A1 (n_3431), .A2 (n_2136));
NOR2_X1 i_1523 (.ZN (n_2531), .A1 (n_3431), .A2 (n_2138));
NOR2_X1 i_1522 (.ZN (n_2530), .A1 (n_3431), .A2 (n_2141));
NOR2_X1 i_1521 (.ZN (n_2529), .A1 (n_3431), .A2 (n_2142));
NOR2_X1 i_1520 (.ZN (n_2528), .A1 (n_3431), .A2 (n_2143));
NOR2_X1 i_1519 (.ZN (n_2527), .A1 (n_3431), .A2 (n_2144));
NOR2_X1 i_1518 (.ZN (n_2526), .A1 (n_3431), .A2 (n_2146));
NOR2_X1 i_1517 (.ZN (n_2525), .A1 (n_3431), .A2 (n_2148));
NOR2_X1 i_1516 (.ZN (n_2523), .A1 (n_3431), .A2 (n_2150));
NOR2_X1 i_1515 (.ZN (n_2521), .A1 (n_3431), .A2 (n_2152));
NOR2_X1 i_1514 (.ZN (n_2520), .A1 (n_3431), .A2 (n_2154));
NOR2_X1 i_1513 (.ZN (n_2519), .A1 (n_3431), .A2 (n_2155));
NOR2_X1 i_1512 (.ZN (n_2518), .A1 (n_3431), .A2 (n_2156));
NOR2_X1 i_1511 (.ZN (n_2517), .A1 (n_3431), .A2 (n_2158));
NOR2_X1 i_1510 (.ZN (n_2516), .A1 (n_3431), .A2 (n_2162));
NOR2_X1 i_1509 (.ZN (n_2515), .A1 (n_3431), .A2 (n_2163));
NOR2_X1 i_1508 (.ZN (n_2514), .A1 (n_3431), .A2 (n_2164));
NOR2_X1 i_1507 (.ZN (n_2513), .A1 (n_3431), .A2 (n_2166));
NOR2_X1 i_1506 (.ZN (n_2512), .A1 (n_3431), .A2 (n_2169));
NOR2_X1 i_1505 (.ZN (n_2511), .A1 (n_3431), .A2 (n_2170));
NOR2_X1 i_1504 (.ZN (n_2510), .A1 (n_3431), .A2 (n_2171));
NOR2_X1 i_1503 (.ZN (n_2509), .A1 (n_3431), .A2 (n_2172));
NOR2_X1 i_1502 (.ZN (n_2508), .A1 (n_3431), .A2 (n_3404));
NOR2_X1 i_1501 (.ZN (n_2507), .A1 (n_3431), .A2 (n_3405));
NOR2_X1 i_1500 (.ZN (n_2506), .A1 (n_3431), .A2 (n_3406));
NOR2_X1 i_1499 (.ZN (n_2505), .A1 (n_3432), .A2 (n_3425));
NOR2_X1 i_1498 (.ZN (n_2504), .A1 (n_3432), .A2 (n_2133));
NOR2_X1 i_1497 (.ZN (n_2503), .A1 (n_3432), .A2 (n_2134));
NOR2_X1 i_1496 (.ZN (n_2502), .A1 (n_3432), .A2 (n_2135));
NOR2_X1 i_1495 (.ZN (n_2501), .A1 (n_3432), .A2 (n_2136));
NOR2_X1 i_1494 (.ZN (n_2500), .A1 (n_3432), .A2 (n_2138));
NOR2_X1 i_1493 (.ZN (n_2499), .A1 (n_3432), .A2 (n_2141));
NOR2_X1 i_1492 (.ZN (n_2498), .A1 (n_3432), .A2 (n_2142));
NOR2_X1 i_1491 (.ZN (n_2497), .A1 (n_3432), .A2 (n_2143));
NOR2_X1 i_1490 (.ZN (n_2496), .A1 (n_3432), .A2 (n_2144));
NOR2_X1 i_1489 (.ZN (n_2495), .A1 (n_3432), .A2 (n_2146));
NOR2_X1 i_1488 (.ZN (n_2493), .A1 (n_3432), .A2 (n_2149));
NOR2_X1 i_1487 (.ZN (n_2491), .A1 (n_3432), .A2 (n_2151));
NOR2_X1 i_1486 (.ZN (n_2490), .A1 (n_3432), .A2 (n_2152));
NOR2_X1 i_1485 (.ZN (n_2489), .A1 (n_3432), .A2 (n_2154));
NOR2_X1 i_1484 (.ZN (n_2488), .A1 (n_3432), .A2 (n_2155));
NOR2_X1 i_1483 (.ZN (n_2487), .A1 (n_3432), .A2 (n_2156));
NOR2_X1 i_1482 (.ZN (n_2486), .A1 (n_3432), .A2 (n_2158));
NOR2_X1 i_1481 (.ZN (n_2485), .A1 (n_3432), .A2 (n_2162));
NOR2_X1 i_1480 (.ZN (n_2484), .A1 (n_3432), .A2 (n_2163));
NOR2_X1 i_1479 (.ZN (n_2483), .A1 (n_3432), .A2 (n_2164));
NOR2_X1 i_1478 (.ZN (n_2482), .A1 (n_3432), .A2 (n_2166));
NOR2_X1 i_1477 (.ZN (n_2481), .A1 (n_3432), .A2 (n_2169));
NOR2_X1 i_1476 (.ZN (n_2480), .A1 (n_3432), .A2 (n_2170));
NOR2_X1 i_1475 (.ZN (n_2479), .A1 (n_3432), .A2 (n_2171));
NOR2_X1 i_1474 (.ZN (n_2478), .A1 (n_3432), .A2 (n_2172));
NOR2_X1 i_1473 (.ZN (n_2477), .A1 (n_3432), .A2 (n_3404));
NOR2_X1 i_1472 (.ZN (n_2476), .A1 (n_3432), .A2 (n_3405));
NOR2_X1 i_1471 (.ZN (n_2475), .A1 (n_3433), .A2 (n_3425));
NOR2_X1 i_1470 (.ZN (n_2474), .A1 (n_3433), .A2 (n_2133));
NOR2_X1 i_1469 (.ZN (n_2473), .A1 (n_3433), .A2 (n_2134));
NOR2_X1 i_1468 (.ZN (n_2472), .A1 (n_3433), .A2 (n_2135));
NOR2_X1 i_1467 (.ZN (n_2471), .A1 (n_3433), .A2 (n_2136));
NOR2_X1 i_1466 (.ZN (n_2470), .A1 (n_3433), .A2 (n_2138));
NOR2_X1 i_1465 (.ZN (n_2469), .A1 (n_3433), .A2 (n_2141));
NOR2_X1 i_1464 (.ZN (n_2468), .A1 (n_3433), .A2 (n_2142));
NOR2_X1 i_1463 (.ZN (n_2467), .A1 (n_3433), .A2 (n_2143));
NOR2_X1 i_1462 (.ZN (n_2466), .A1 (n_3433), .A2 (n_2144));
NOR2_X1 i_1461 (.ZN (n_2464), .A1 (n_3433), .A2 (n_2148));
NOR2_X1 i_1460 (.ZN (n_2462), .A1 (n_3433), .A2 (n_2150));
NOR2_X1 i_1459 (.ZN (n_2461), .A1 (n_3433), .A2 (n_2151));
NOR2_X1 i_1458 (.ZN (n_2460), .A1 (n_3433), .A2 (n_2152));
NOR2_X1 i_1457 (.ZN (n_2459), .A1 (n_3433), .A2 (n_2154));
NOR2_X1 i_1456 (.ZN (n_2458), .A1 (n_3433), .A2 (n_2155));
NOR2_X1 i_1455 (.ZN (n_2457), .A1 (n_3433), .A2 (n_2156));
NOR2_X1 i_1454 (.ZN (n_2456), .A1 (n_3433), .A2 (n_2158));
NOR2_X1 i_1453 (.ZN (n_2455), .A1 (n_3433), .A2 (n_2162));
NOR2_X1 i_1452 (.ZN (n_2454), .A1 (n_3433), .A2 (n_2163));
NOR2_X1 i_1451 (.ZN (n_2453), .A1 (n_3433), .A2 (n_2164));
NOR2_X1 i_1450 (.ZN (n_2452), .A1 (n_3433), .A2 (n_2166));
NOR2_X1 i_1449 (.ZN (n_2451), .A1 (n_3433), .A2 (n_2169));
NOR2_X1 i_1448 (.ZN (n_2450), .A1 (n_3433), .A2 (n_2170));
NOR2_X1 i_1447 (.ZN (n_2449), .A1 (n_3433), .A2 (n_2171));
NOR2_X1 i_1446 (.ZN (n_2448), .A1 (n_3433), .A2 (n_2172));
NOR2_X1 i_1445 (.ZN (n_2447), .A1 (n_3433), .A2 (n_3404));
NOR2_X1 i_1444 (.ZN (n_2446), .A1 (n_3434), .A2 (n_3425));
NOR2_X1 i_1443 (.ZN (n_2445), .A1 (n_3434), .A2 (n_2133));
NOR2_X1 i_1442 (.ZN (n_2444), .A1 (n_3434), .A2 (n_2134));
NOR2_X1 i_1441 (.ZN (n_2443), .A1 (n_3434), .A2 (n_2135));
NOR2_X1 i_1440 (.ZN (n_2442), .A1 (n_3434), .A2 (n_2136));
NOR2_X1 i_1439 (.ZN (n_2441), .A1 (n_3434), .A2 (n_2138));
NOR2_X1 i_1438 (.ZN (n_2440), .A1 (n_3434), .A2 (n_2141));
NOR2_X1 i_1437 (.ZN (n_2439), .A1 (n_3434), .A2 (n_2142));
NOR2_X1 i_1436 (.ZN (n_2438), .A1 (n_3434), .A2 (n_2143));
NOR2_X1 i_1435 (.ZN (n_2436), .A1 (n_3434), .A2 (n_2146));
NOR2_X1 i_1434 (.ZN (n_2434), .A1 (n_3434), .A2 (n_2149));
NOR2_X1 i_1433 (.ZN (n_2433), .A1 (n_3434), .A2 (n_2150));
NOR2_X1 i_1432 (.ZN (n_2432), .A1 (n_3434), .A2 (n_2151));
NOR2_X1 i_1431 (.ZN (n_2431), .A1 (n_3434), .A2 (n_2152));
NOR2_X1 i_1430 (.ZN (n_2430), .A1 (n_3434), .A2 (n_2154));
NOR2_X1 i_1429 (.ZN (n_2429), .A1 (n_3434), .A2 (n_2155));
NOR2_X1 i_1428 (.ZN (n_2428), .A1 (n_3434), .A2 (n_2156));
NOR2_X1 i_1427 (.ZN (n_2427), .A1 (n_3434), .A2 (n_2158));
NOR2_X1 i_1426 (.ZN (n_2426), .A1 (n_3434), .A2 (n_2162));
NOR2_X1 i_1425 (.ZN (n_2425), .A1 (n_3434), .A2 (n_2163));
NOR2_X1 i_1424 (.ZN (n_2424), .A1 (n_3434), .A2 (n_2164));
NOR2_X1 i_1423 (.ZN (n_2423), .A1 (n_3434), .A2 (n_2166));
NOR2_X1 i_1422 (.ZN (n_2422), .A1 (n_3434), .A2 (n_2169));
NOR2_X1 i_1421 (.ZN (n_2421), .A1 (n_3434), .A2 (n_2170));
NOR2_X1 i_1420 (.ZN (n_2420), .A1 (n_3434), .A2 (n_2171));
NOR2_X1 i_1419 (.ZN (n_2419), .A1 (n_3434), .A2 (n_2172));
NOR2_X1 i_1418 (.ZN (n_2418), .A1 (n_3434), .A2 (n_3404));
NOR2_X1 i_1417 (.ZN (n_2417), .A1 (n_3434), .A2 (n_3405));
NOR2_X1 i_1416 (.ZN (n_2416), .A1 (n_3434), .A2 (n_3406));
NOR2_X1 i_1415 (.ZN (n_2415), .A1 (n_3435), .A2 (n_3425));
NOR2_X1 i_1414 (.ZN (n_2414), .A1 (n_3435), .A2 (n_2133));
NOR2_X1 i_1413 (.ZN (n_2413), .A1 (n_3435), .A2 (n_2134));
NOR2_X1 i_1412 (.ZN (n_2412), .A1 (n_3435), .A2 (n_2135));
NOR2_X1 i_1411 (.ZN (n_2411), .A1 (n_3435), .A2 (n_2136));
NOR2_X1 i_1410 (.ZN (n_2410), .A1 (n_3435), .A2 (n_2138));
NOR2_X1 i_1409 (.ZN (n_2409), .A1 (n_3435), .A2 (n_2141));
NOR2_X1 i_1408 (.ZN (n_2408), .A1 (n_3435), .A2 (n_2142));
NOR2_X1 i_1407 (.ZN (n_2406), .A1 (n_3435), .A2 (n_2144));
NOR2_X1 i_1406 (.ZN (n_2404), .A1 (n_3435), .A2 (n_2148));
NOR2_X1 i_1405 (.ZN (n_2403), .A1 (n_3435), .A2 (n_2149));
NOR2_X1 i_1404 (.ZN (n_2402), .A1 (n_3435), .A2 (n_2150));
NOR2_X1 i_1403 (.ZN (n_2401), .A1 (n_3435), .A2 (n_2151));
NOR2_X1 i_1402 (.ZN (n_2400), .A1 (n_3435), .A2 (n_2152));
NOR2_X1 i_1401 (.ZN (n_2399), .A1 (n_3435), .A2 (n_2154));
NOR2_X1 i_1400 (.ZN (n_2398), .A1 (n_3435), .A2 (n_2155));
NOR2_X1 i_1399 (.ZN (n_2397), .A1 (n_3435), .A2 (n_2156));
NOR2_X1 i_1398 (.ZN (n_2396), .A1 (n_3435), .A2 (n_2158));
NOR2_X1 i_1397 (.ZN (n_2395), .A1 (n_3435), .A2 (n_2162));
NOR2_X1 i_1396 (.ZN (n_2394), .A1 (n_3435), .A2 (n_2163));
NOR2_X1 i_1395 (.ZN (n_2393), .A1 (n_3435), .A2 (n_2164));
NOR2_X1 i_1394 (.ZN (n_2392), .A1 (n_3435), .A2 (n_2166));
NOR2_X1 i_1393 (.ZN (n_2391), .A1 (n_3435), .A2 (n_2169));
NOR2_X1 i_1392 (.ZN (n_2390), .A1 (n_3435), .A2 (n_2170));
NOR2_X1 i_1391 (.ZN (n_2389), .A1 (n_3435), .A2 (n_2171));
NOR2_X1 i_1390 (.ZN (n_2388), .A1 (n_3435), .A2 (n_2172));
NOR2_X1 i_1389 (.ZN (n_2387), .A1 (n_3435), .A2 (n_3404));
NOR2_X1 i_1388 (.ZN (n_2386), .A1 (n_3435), .A2 (n_3405));
NOR2_X1 i_1387 (.ZN (n_2385), .A1 (n_3436), .A2 (n_3425));
NOR2_X1 i_1386 (.ZN (n_2384), .A1 (n_3436), .A2 (n_2133));
NOR2_X1 i_1385 (.ZN (n_2383), .A1 (n_3436), .A2 (n_2134));
NOR2_X1 i_1384 (.ZN (n_2382), .A1 (n_3436), .A2 (n_2135));
NOR2_X1 i_1383 (.ZN (n_2381), .A1 (n_3436), .A2 (n_2136));
NOR2_X1 i_1382 (.ZN (n_2380), .A1 (n_3436), .A2 (n_2138));
NOR2_X1 i_1381 (.ZN (n_2379), .A1 (n_3436), .A2 (n_2141));
NOR2_X1 i_1380 (.ZN (n_2377), .A1 (n_3436), .A2 (n_2143));
NOR2_X1 i_1379 (.ZN (n_2375), .A1 (n_3436), .A2 (n_2146));
NOR2_X1 i_1378 (.ZN (n_2374), .A1 (n_3436), .A2 (n_2148));
NOR2_X1 i_1377 (.ZN (n_2373), .A1 (n_3436), .A2 (n_2149));
NOR2_X1 i_1376 (.ZN (n_2372), .A1 (n_3436), .A2 (n_2150));
NOR2_X1 i_1375 (.ZN (n_2371), .A1 (n_3436), .A2 (n_2151));
NOR2_X1 i_1374 (.ZN (n_2370), .A1 (n_3436), .A2 (n_2152));
NOR2_X1 i_1373 (.ZN (n_2369), .A1 (n_3436), .A2 (n_2154));
NOR2_X1 i_1372 (.ZN (n_2368), .A1 (n_3436), .A2 (n_2155));
NOR2_X1 i_1371 (.ZN (n_2367), .A1 (n_3436), .A2 (n_2156));
NOR2_X1 i_1370 (.ZN (n_2366), .A1 (n_3436), .A2 (n_2158));
NOR2_X1 i_1369 (.ZN (n_2365), .A1 (n_3436), .A2 (n_2162));
NOR2_X1 i_1368 (.ZN (n_2364), .A1 (n_3436), .A2 (n_2163));
NOR2_X1 i_1367 (.ZN (n_2363), .A1 (n_3436), .A2 (n_2164));
NOR2_X1 i_1366 (.ZN (n_2362), .A1 (n_3436), .A2 (n_2166));
NOR2_X1 i_1365 (.ZN (n_2361), .A1 (n_3436), .A2 (n_2169));
NOR2_X1 i_1364 (.ZN (n_2360), .A1 (n_3436), .A2 (n_2170));
NOR2_X1 i_1363 (.ZN (n_2359), .A1 (n_3436), .A2 (n_2171));
NOR2_X1 i_1362 (.ZN (n_2358), .A1 (n_3436), .A2 (n_2172));
NOR2_X1 i_1361 (.ZN (n_2357), .A1 (n_3436), .A2 (n_3404));
NOR2_X1 i_1360 (.ZN (n_2356), .A1 (n_3437), .A2 (n_3425));
NOR2_X1 i_1359 (.ZN (n_2355), .A1 (n_3437), .A2 (n_2133));
NOR2_X1 i_1358 (.ZN (n_2354), .A1 (n_3437), .A2 (n_2134));
NOR2_X1 i_1357 (.ZN (n_2353), .A1 (n_3437), .A2 (n_2135));
NOR2_X1 i_1356 (.ZN (n_2352), .A1 (n_3437), .A2 (n_2136));
NOR2_X1 i_1355 (.ZN (n_2351), .A1 (n_3437), .A2 (n_2138));
NOR2_X1 i_1354 (.ZN (n_2349), .A1 (n_3437), .A2 (n_2142));
NOR2_X1 i_1353 (.ZN (n_2347), .A1 (n_3437), .A2 (n_2144));
NOR2_X1 i_1352 (.ZN (n_2345), .A1 (n_3437), .A2 (n_2148));
NOR2_X1 i_1351 (.ZN (n_2344), .A1 (n_3437), .A2 (n_2149));
NOR2_X1 i_1350 (.ZN (n_2343), .A1 (n_3437), .A2 (n_2150));
NOR2_X1 i_1349 (.ZN (n_2342), .A1 (n_3437), .A2 (n_2151));
NOR2_X1 i_1348 (.ZN (n_2341), .A1 (n_3437), .A2 (n_2152));
NOR2_X1 i_1347 (.ZN (n_2340), .A1 (n_3437), .A2 (n_2154));
NOR2_X1 i_1346 (.ZN (n_2339), .A1 (n_3437), .A2 (n_2155));
NOR2_X1 i_1345 (.ZN (n_2338), .A1 (n_3437), .A2 (n_2156));
NOR2_X1 i_1344 (.ZN (n_2337), .A1 (n_3437), .A2 (n_2158));
NOR2_X1 i_1343 (.ZN (n_2336), .A1 (n_3437), .A2 (n_2162));
NOR2_X1 i_1342 (.ZN (n_2335), .A1 (n_3437), .A2 (n_2163));
NOR2_X1 i_1341 (.ZN (n_2334), .A1 (n_3437), .A2 (n_2164));
NOR2_X1 i_1340 (.ZN (n_2333), .A1 (n_3437), .A2 (n_2166));
NOR2_X1 i_1339 (.ZN (n_2332), .A1 (n_3437), .A2 (n_2169));
NOR2_X1 i_1338 (.ZN (n_2331), .A1 (n_3437), .A2 (n_2170));
NOR2_X1 i_1337 (.ZN (n_2330), .A1 (n_3437), .A2 (n_2171));
NOR2_X1 i_1336 (.ZN (n_2329), .A1 (n_3437), .A2 (n_2172));
NOR2_X1 i_1335 (.ZN (n_2328), .A1 (n_3437), .A2 (n_3404));
NOR2_X1 i_1334 (.ZN (n_2327), .A1 (n_3437), .A2 (n_3405));
NOR2_X1 i_1333 (.ZN (n_2326), .A1 (n_3437), .A2 (n_3406));
NOR2_X1 i_1332 (.ZN (n_2325), .A1 (n_3438), .A2 (n_3425));
NOR2_X1 i_1331 (.ZN (n_2324), .A1 (n_3438), .A2 (n_2133));
NOR2_X1 i_1330 (.ZN (n_2323), .A1 (n_3438), .A2 (n_2134));
NOR2_X1 i_1329 (.ZN (n_2322), .A1 (n_3438), .A2 (n_2135));
NOR2_X1 i_1328 (.ZN (n_2321), .A1 (n_3438), .A2 (n_2136));
NOR2_X1 i_1327 (.ZN (n_2320), .A1 (n_3438), .A2 (n_2138));
NOR2_X1 i_1326 (.ZN (n_2319), .A1 (n_3438), .A2 (n_2141));
NOR2_X1 i_1325 (.ZN (n_2317), .A1 (n_3438), .A2 (n_2143));
NOR2_X1 i_1324 (.ZN (n_2315), .A1 (n_3438), .A2 (n_2146));
NOR2_X1 i_1323 (.ZN (n_2314), .A1 (n_3438), .A2 (n_2148));
NOR2_X1 i_1322 (.ZN (n_2313), .A1 (n_3438), .A2 (n_2149));
NOR2_X1 i_1321 (.ZN (n_2312), .A1 (n_3438), .A2 (n_2150));
NOR2_X1 i_1320 (.ZN (n_2311), .A1 (n_3438), .A2 (n_2151));
NOR2_X1 i_1319 (.ZN (n_2310), .A1 (n_3438), .A2 (n_2152));
NOR2_X1 i_1318 (.ZN (n_2309), .A1 (n_3438), .A2 (n_2154));
NOR2_X1 i_1317 (.ZN (n_2308), .A1 (n_3438), .A2 (n_2155));
NOR2_X1 i_1316 (.ZN (n_2307), .A1 (n_3438), .A2 (n_2156));
NOR2_X1 i_1315 (.ZN (n_2306), .A1 (n_3438), .A2 (n_2158));
NOR2_X1 i_1314 (.ZN (n_2305), .A1 (n_3438), .A2 (n_2162));
NOR2_X1 i_1313 (.ZN (n_2304), .A1 (n_3438), .A2 (n_2163));
NOR2_X1 i_1312 (.ZN (n_2303), .A1 (n_3438), .A2 (n_2164));
NOR2_X1 i_1311 (.ZN (n_2302), .A1 (n_3438), .A2 (n_2166));
NOR2_X1 i_1310 (.ZN (n_2301), .A1 (n_3438), .A2 (n_2169));
NOR2_X1 i_1309 (.ZN (n_2300), .A1 (n_3438), .A2 (n_2170));
NOR2_X1 i_1308 (.ZN (n_2299), .A1 (n_3438), .A2 (n_2171));
NOR2_X1 i_1307 (.ZN (n_2298), .A1 (n_3438), .A2 (n_2172));
NOR2_X1 i_1306 (.ZN (n_2297), .A1 (n_3438), .A2 (n_3404));
NOR2_X1 i_1305 (.ZN (n_2296), .A1 (n_3438), .A2 (n_3405));
NOR2_X1 i_1304 (.ZN (n_2295), .A1 (n_3439), .A2 (n_3425));
NOR2_X1 i_1303 (.ZN (n_2294), .A1 (n_3439), .A2 (n_2133));
NOR2_X1 i_1302 (.ZN (n_2293), .A1 (n_3439), .A2 (n_2134));
NOR2_X1 i_1301 (.ZN (n_2292), .A1 (n_3439), .A2 (n_2135));
NOR2_X1 i_1300 (.ZN (n_2291), .A1 (n_3439), .A2 (n_2136));
NOR2_X1 i_1299 (.ZN (n_2290), .A1 (n_3439), .A2 (n_2138));
NOR2_X1 i_1298 (.ZN (n_2288), .A1 (n_3439), .A2 (n_2142));
NOR2_X1 i_1297 (.ZN (n_2286), .A1 (n_3439), .A2 (n_2144));
NOR2_X1 i_1296 (.ZN (n_2285), .A1 (n_3439), .A2 (n_2146));
NOR2_X1 i_1295 (.ZN (n_2284), .A1 (n_3439), .A2 (n_2148));
NOR2_X1 i_1294 (.ZN (n_2283), .A1 (n_3439), .A2 (n_2149));
NOR2_X1 i_1293 (.ZN (n_2282), .A1 (n_3439), .A2 (n_2150));
NOR2_X1 i_1292 (.ZN (n_2281), .A1 (n_3439), .A2 (n_2151));
NOR2_X1 i_1291 (.ZN (n_2280), .A1 (n_3439), .A2 (n_2152));
NOR2_X1 i_1290 (.ZN (n_2279), .A1 (n_3439), .A2 (n_2154));
NOR2_X1 i_1289 (.ZN (n_2278), .A1 (n_3439), .A2 (n_2155));
NOR2_X1 i_1288 (.ZN (n_2277), .A1 (n_3439), .A2 (n_2156));
NOR2_X1 i_1287 (.ZN (n_2276), .A1 (n_3439), .A2 (n_2158));
NOR2_X1 i_1286 (.ZN (n_2275), .A1 (n_3439), .A2 (n_2162));
NOR2_X1 i_1285 (.ZN (n_2274), .A1 (n_3439), .A2 (n_2163));
NOR2_X1 i_1284 (.ZN (n_2273), .A1 (n_3439), .A2 (n_2164));
NOR2_X1 i_1283 (.ZN (n_2272), .A1 (n_3439), .A2 (n_2166));
NOR2_X1 i_1282 (.ZN (n_2271), .A1 (n_3439), .A2 (n_2169));
NOR2_X1 i_1281 (.ZN (n_2270), .A1 (n_3439), .A2 (n_2170));
NOR2_X1 i_1280 (.ZN (n_2269), .A1 (n_3439), .A2 (n_2171));
NOR2_X1 i_1279 (.ZN (n_2268), .A1 (n_3439), .A2 (n_2172));
NOR2_X1 i_1278 (.ZN (n_2267), .A1 (n_3439), .A2 (n_3404));
NOR2_X1 i_1277 (.ZN (n_2266), .A1 (n_3440), .A2 (n_3425));
NOR2_X1 i_1276 (.ZN (n_2265), .A1 (n_3440), .A2 (n_2133));
NOR2_X1 i_1275 (.ZN (n_2264), .A1 (n_3440), .A2 (n_2134));
NOR2_X1 i_1274 (.ZN (n_2263), .A1 (n_3440), .A2 (n_2135));
NOR2_X1 i_1273 (.ZN (n_2262), .A1 (n_3440), .A2 (n_2136));
NOR2_X1 i_1272 (.ZN (n_2260), .A1 (n_3440), .A2 (n_2141));
NOR2_X1 i_1271 (.ZN (n_2258), .A1 (n_3440), .A2 (n_2143));
NOR2_X1 i_1270 (.ZN (n_2257), .A1 (n_3440), .A2 (n_2144));
NOR2_X1 i_1269 (.ZN (n_2256), .A1 (n_3440), .A2 (n_2146));
NOR2_X1 i_1268 (.ZN (n_2255), .A1 (n_3440), .A2 (n_2148));
NOR2_X1 i_1267 (.ZN (n_2254), .A1 (n_3440), .A2 (n_2149));
NOR2_X1 i_1266 (.ZN (n_2253), .A1 (n_3440), .A2 (n_2150));
NOR2_X1 i_1265 (.ZN (n_2252), .A1 (n_3440), .A2 (n_2151));
NOR2_X1 i_1264 (.ZN (n_2251), .A1 (n_3440), .A2 (n_2152));
NOR2_X1 i_1263 (.ZN (n_2250), .A1 (n_3440), .A2 (n_2154));
NOR2_X1 i_1262 (.ZN (n_2249), .A1 (n_3440), .A2 (n_2155));
NOR2_X1 i_1261 (.ZN (n_2248), .A1 (n_3440), .A2 (n_2156));
NOR2_X1 i_1260 (.ZN (n_2247), .A1 (n_3440), .A2 (n_2158));
NOR2_X1 i_1259 (.ZN (n_2246), .A1 (n_3440), .A2 (n_2162));
NOR2_X1 i_1258 (.ZN (n_2245), .A1 (n_3440), .A2 (n_2163));
NOR2_X1 i_1257 (.ZN (n_2244), .A1 (n_3440), .A2 (n_2164));
NOR2_X1 i_1256 (.ZN (n_2243), .A1 (n_3440), .A2 (n_2166));
NOR2_X1 i_1255 (.ZN (n_2242), .A1 (n_3440), .A2 (n_2169));
NOR2_X1 i_1254 (.ZN (n_2241), .A1 (n_3440), .A2 (n_2170));
NOR2_X1 i_1253 (.ZN (n_2240), .A1 (n_3440), .A2 (n_2171));
NOR2_X1 i_1252 (.ZN (n_2239), .A1 (n_3440), .A2 (n_2172));
NOR2_X1 i_1251 (.ZN (n_2238), .A1 (n_3440), .A2 (n_3404));
NOR2_X1 i_1250 (.ZN (n_2237), .A1 (n_3440), .A2 (n_3405));
NOR2_X1 i_1249 (.ZN (n_2236), .A1 (n_3440), .A2 (n_3406));
NOR2_X1 i_1248 (.ZN (n_2235), .A1 (n_3441), .A2 (n_3425));
NOR2_X1 i_1247 (.ZN (n_2234), .A1 (n_3441), .A2 (n_2133));
NOR2_X1 i_1246 (.ZN (n_2233), .A1 (n_3441), .A2 (n_2134));
NOR2_X1 i_1245 (.ZN (n_2232), .A1 (n_3441), .A2 (n_2135));
NOR2_X1 i_1244 (.ZN (n_2230), .A1 (n_3441), .A2 (n_2138));
NOR2_X1 i_1243 (.ZN (n_2228), .A1 (n_3441), .A2 (n_2142));
NOR2_X1 i_1242 (.ZN (n_2227), .A1 (n_3441), .A2 (n_2143));
NOR2_X1 i_1241 (.ZN (n_2226), .A1 (n_3441), .A2 (n_2144));
NOR2_X1 i_1240 (.ZN (n_2225), .A1 (n_3441), .A2 (n_2146));
NOR2_X1 i_1239 (.ZN (n_2224), .A1 (n_3441), .A2 (n_2148));
NOR2_X1 i_1238 (.ZN (n_2223), .A1 (n_3441), .A2 (n_2149));
NOR2_X1 i_1237 (.ZN (n_2222), .A1 (n_3441), .A2 (n_2150));
NOR2_X1 i_1236 (.ZN (n_2221), .A1 (n_3441), .A2 (n_2151));
NOR2_X1 i_1235 (.ZN (n_2220), .A1 (n_3441), .A2 (n_2152));
NOR2_X1 i_1234 (.ZN (n_2219), .A1 (n_3441), .A2 (n_2154));
NOR2_X1 i_1233 (.ZN (n_2218), .A1 (n_3441), .A2 (n_2155));
NOR2_X1 i_1232 (.ZN (n_2217), .A1 (n_3441), .A2 (n_2156));
NOR2_X1 i_1231 (.ZN (n_2216), .A1 (n_3441), .A2 (n_2158));
NOR2_X1 i_1230 (.ZN (n_2215), .A1 (n_3441), .A2 (n_2162));
NOR2_X1 i_1229 (.ZN (n_2214), .A1 (n_3441), .A2 (n_2163));
NOR2_X1 i_1228 (.ZN (n_2213), .A1 (n_3441), .A2 (n_2164));
NOR2_X1 i_1227 (.ZN (n_2212), .A1 (n_3441), .A2 (n_2166));
NOR2_X1 i_1226 (.ZN (n_2211), .A1 (n_3441), .A2 (n_2169));
NOR2_X1 i_1225 (.ZN (n_2210), .A1 (n_3441), .A2 (n_2170));
NOR2_X1 i_1224 (.ZN (n_2209), .A1 (n_3441), .A2 (n_2171));
NOR2_X1 i_1223 (.ZN (n_2208), .A1 (n_3441), .A2 (n_2172));
NOR2_X1 i_1222 (.ZN (n_2207), .A1 (n_3441), .A2 (n_3404));
NOR2_X1 i_1221 (.ZN (n_2206), .A1 (n_3441), .A2 (n_3405));
NOR2_X1 i_1220 (.ZN (n_2205), .A1 (n_3442), .A2 (n_3425));
NOR2_X1 i_1219 (.ZN (n_2204), .A1 (n_3442), .A2 (n_2133));
NOR2_X1 i_1218 (.ZN (n_2203), .A1 (n_3442), .A2 (n_2134));
NOR2_X1 i_1217 (.ZN (n_2201), .A1 (n_3442), .A2 (n_2136));
NOR2_X1 i_1216 (.ZN (n_2199), .A1 (n_3442), .A2 (n_2141));
NOR2_X1 i_1215 (.ZN (n_2198), .A1 (n_3442), .A2 (n_2142));
NOR2_X1 i_1214 (.ZN (n_2197), .A1 (n_3442), .A2 (n_2143));
NOR2_X1 i_1213 (.ZN (n_2196), .A1 (n_3442), .A2 (n_2144));
NOR2_X1 i_1212 (.ZN (n_2195), .A1 (n_3442), .A2 (n_2146));
NOR2_X1 i_1211 (.ZN (n_2194), .A1 (n_3442), .A2 (n_2148));
NOR2_X1 i_1210 (.ZN (n_2193), .A1 (n_3442), .A2 (n_2149));
NOR2_X1 i_1209 (.ZN (n_2192), .A1 (n_3442), .A2 (n_2150));
NOR2_X1 i_1208 (.ZN (n_2191), .A1 (n_3442), .A2 (n_2151));
NOR2_X1 i_1207 (.ZN (n_2190), .A1 (n_3442), .A2 (n_2152));
NOR2_X1 i_1206 (.ZN (n_2189), .A1 (n_3442), .A2 (n_2154));
NOR2_X1 i_1205 (.ZN (n_2188), .A1 (n_3442), .A2 (n_2155));
NOR2_X1 i_1204 (.ZN (n_2187), .A1 (n_3442), .A2 (n_2156));
NOR2_X1 i_1203 (.ZN (n_2186), .A1 (n_3442), .A2 (n_2158));
NOR2_X1 i_1202 (.ZN (n_2185), .A1 (n_3442), .A2 (n_2162));
NOR2_X1 i_1201 (.ZN (n_2184), .A1 (n_3442), .A2 (n_2163));
NOR2_X1 i_1200 (.ZN (n_2183), .A1 (n_3442), .A2 (n_2164));
NOR2_X1 i_1199 (.ZN (n_2182), .A1 (n_3442), .A2 (n_2166));
NOR2_X1 i_1198 (.ZN (n_2181), .A1 (n_3442), .A2 (n_2169));
NOR2_X1 i_1197 (.ZN (n_2180), .A1 (n_3442), .A2 (n_2170));
NOR2_X1 i_1196 (.ZN (n_2179), .A1 (n_3442), .A2 (n_2171));
NOR2_X1 i_1195 (.ZN (n_2178), .A1 (n_3442), .A2 (n_2172));
NOR2_X1 i_1194 (.ZN (n_2177), .A1 (n_3442), .A2 (n_3404));
NOR2_X1 i_1193 (.ZN (n_2176), .A1 (n_3443), .A2 (n_3425));
NOR2_X1 i_1192 (.ZN (n_2175), .A1 (n_3443), .A2 (n_2133));
NOR2_X1 i_1191 (.ZN (n_2174), .A1 (n_3443), .A2 (n_2135));
NOR2_X1 i_1190 (.ZN (n_2173), .A1 (n_3444), .A2 (n_3425));
OAI21_X1 i_1189 (.ZN (n_2168), .A (n_1773), .B1 (n_1776), .B2 (n_1775));
XNOR2_X1 i_1188 (.ZN (n_2167), .A (n_1772), .B (n_2168));
INV_X1 i_1187 (.ZN (n_2161), .A (n_1766));
NOR2_X1 i_1186 (.ZN (n_2160), .A1 (n_1763), .A2 (n_2161));
XOR2_X1 i_1185 (.Z (n_2159), .A (n_984), .B (n_2160));
OAI21_X1 i_1184 (.ZN (n_2153), .A (n_1777), .B1 (n_2126), .B2 (n_2125));
OAI21_X1 i_1183 (.ZN (n_2140), .A (n_1768), .B1 (n_1770), .B2 (n_1769));
XNOR2_X1 i_1182 (.ZN (n_2139), .A (n_1767), .B (n_2140));
NOR2_X1 i_1181 (.ZN (n_2131), .A1 (n_1759), .A2 (n_1757));
OAI21_X1 i_1180 (.ZN (n_2123), .A (n_2132), .B1 (n_2129), .B2 (n_2128));
NAND2_X1 i_1179 (.ZN (n_2122), .A1 (n_2127), .A2 (n_2123));
NOR2_X1 i_1178 (.ZN (n_2121), .A1 (n_3414), .A2 (n_3410));
NAND2_X1 i_1177 (.ZN (n_2120), .A1 (n_1762), .A2 (n_2121));
INV_X1 i_1176 (.ZN (n_2119), .A (n_2120));
OAI21_X1 i_1175 (.ZN (n_2118), .A (n_2120), .B1 (n_1762), .B2 (n_2121));
NOR2_X1 i_1174 (.ZN (n_2117), .A1 (n_1761), .A2 (n_2131));
XOR2_X1 i_1173 (.Z (n_2116), .A (n_2118), .B (n_2117));
OAI22_X1 i_1172 (.ZN (n_2115), .A1 (n_1762), .A2 (n_2121), .B1 (n_2119), .B2 (n_2117));
NOR2_X1 i_1171 (.ZN (n_2114), .A1 (n_3443), .A2 (n_2141));
NAND2_X1 i_1170 (.ZN (n_2113), .A1 (inputB[31]), .A2 (inputA[4]));
NOR2_X1 i_1169 (.ZN (n_2112), .A1 (n_3444), .A2 (n_2138));
NAND2_X1 i_1168 (.ZN (n_2111), .A1 (n_2113), .A2 (n_2112));
OAI21_X1 i_1167 (.ZN (n_2110), .A (n_2111), .B1 (n_2113), .B2 (n_2112));
XNOR2_X1 i_1166 (.ZN (n_2109), .A (n_2114), .B (n_2110));
OAI21_X1 i_1165 (.ZN (n_2108), .A (n_2114), .B1 (n_2113), .B2 (n_2112));
NAND2_X1 i_1164 (.ZN (n_2107), .A1 (n_2111), .A2 (n_2108));
NAND2_X1 i_1163 (.ZN (n_2106), .A1 (inputB[4]), .A2 (inputA[31]));
AND2_X1 i_1162 (.ZN (n_2105), .A1 (n_1049), .A2 (n_2106));
NOR2_X1 i_1161 (.ZN (n_2104), .A1 (n_1049), .A2 (n_2106));
NOR2_X1 i_1160 (.ZN (n_2103), .A1 (n_2105), .A2 (n_2104));
XOR2_X1 i_1159 (.Z (n_2102), .A (n_1051), .B (n_2103));
NOR2_X1 i_1158 (.ZN (n_2101), .A1 (n_1051), .A2 (n_2105));
NOR2_X1 i_1157 (.ZN (n_2100), .A1 (n_2104), .A2 (n_2101));
NOR2_X1 i_1156 (.ZN (n_2099), .A1 (n_3443), .A2 (n_2142));
NAND2_X1 i_1155 (.ZN (n_2098), .A1 (inputB[31]), .A2 (inputA[5]));
NOR2_X1 i_1154 (.ZN (n_2097), .A1 (n_3444), .A2 (n_2141));
NAND2_X1 i_1153 (.ZN (n_2096), .A1 (n_2098), .A2 (n_2097));
OAI21_X1 i_1152 (.ZN (n_2095), .A (n_2096), .B1 (n_2098), .B2 (n_2097));
XNOR2_X1 i_1151 (.ZN (n_2094), .A (n_2099), .B (n_2095));
OAI21_X1 i_1150 (.ZN (n_2093), .A (n_2099), .B1 (n_2098), .B2 (n_2097));
NAND2_X1 i_1149 (.ZN (n_2092), .A1 (n_2096), .A2 (n_2093));
NAND2_X1 i_1148 (.ZN (n_2091), .A1 (inputB[7]), .A2 (inputA[30]));
NOR3_X1 i_1147 (.ZN (n_2090), .A1 (n_3417), .A2 (n_3405), .A3 (n_2091));
AOI22_X1 i_1146 (.ZN (n_2089), .A1 (inputB[7]), .A2 (inputA[29]), .B1 (inputB[6]), .B2 (inputA[30]));
NOR2_X1 i_1145 (.ZN (n_2088), .A1 (n_2090), .A2 (n_2089));
NOR2_X1 i_1144 (.ZN (n_2087), .A1 (n_3416), .A2 (n_3410));
NOR2_X1 i_1143 (.ZN (n_2086), .A1 (n_2089), .A2 (n_2087));
XNOR2_X1 i_1142 (.ZN (n_2085), .A (n_2088), .B (n_2087));
NOR2_X1 i_1141 (.ZN (n_2084), .A1 (n_3443), .A2 (n_2143));
NAND2_X1 i_1140 (.ZN (n_2083), .A1 (inputB[31]), .A2 (inputA[6]));
NOR2_X1 i_1139 (.ZN (n_2082), .A1 (n_3444), .A2 (n_2142));
NAND2_X1 i_1138 (.ZN (n_2081), .A1 (n_2083), .A2 (n_2082));
OAI21_X1 i_1137 (.ZN (n_2080), .A (n_2081), .B1 (n_2083), .B2 (n_2082));
XNOR2_X1 i_1136 (.ZN (n_2079), .A (n_2084), .B (n_2080));
OAI21_X1 i_1135 (.ZN (n_2078), .A (n_2084), .B1 (n_2083), .B2 (n_2082));
NAND2_X1 i_1134 (.ZN (n_2077), .A1 (n_2081), .A2 (n_2078));
NOR2_X1 i_1133 (.ZN (n_2076), .A1 (n_3417), .A2 (n_3410));
NAND2_X1 i_1132 (.ZN (n_2075), .A1 (n_2091), .A2 (n_2076));
INV_X1 i_1131 (.ZN (n_2074), .A (n_2075));
OAI21_X1 i_1130 (.ZN (n_2073), .A (n_2075), .B1 (n_2091), .B2 (n_2076));
NOR2_X1 i_1129 (.ZN (n_2072), .A1 (n_2090), .A2 (n_2086));
XOR2_X1 i_1128 (.Z (n_2071), .A (n_2073), .B (n_2072));
OAI22_X1 i_1127 (.ZN (n_2070), .A1 (n_2091), .A2 (n_2076), .B1 (n_2074), .B2 (n_2072));
NOR2_X1 i_1126 (.ZN (n_2069), .A1 (n_3443), .A2 (n_2144));
NAND2_X1 i_1125 (.ZN (n_2068), .A1 (inputB[31]), .A2 (inputA[7]));
NOR2_X1 i_1124 (.ZN (n_2067), .A1 (n_3444), .A2 (n_2143));
NAND2_X1 i_1123 (.ZN (n_2066), .A1 (n_2068), .A2 (n_2067));
OAI21_X1 i_1122 (.ZN (n_2065), .A (n_2066), .B1 (n_2068), .B2 (n_2067));
XNOR2_X1 i_1121 (.ZN (n_2064), .A (n_2069), .B (n_2065));
OAI21_X1 i_1120 (.ZN (n_2063), .A (n_2069), .B1 (n_2068), .B2 (n_2067));
NAND2_X1 i_1119 (.ZN (n_2062), .A1 (n_2066), .A2 (n_2063));
NAND2_X1 i_1118 (.ZN (n_2061), .A1 (inputB[7]), .A2 (inputA[31]));
AND2_X1 i_1117 (.ZN (n_2060), .A1 (n_1197), .A2 (n_2061));
NOR2_X1 i_1116 (.ZN (n_2059), .A1 (n_1197), .A2 (n_2061));
NOR2_X1 i_1115 (.ZN (n_2058), .A1 (n_2060), .A2 (n_2059));
XOR2_X1 i_1114 (.Z (n_2057), .A (n_1199), .B (n_2058));
NOR2_X1 i_1113 (.ZN (n_2056), .A1 (n_1199), .A2 (n_2060));
NOR2_X1 i_1112 (.ZN (n_2055), .A1 (n_2059), .A2 (n_2056));
NOR2_X1 i_1111 (.ZN (n_2054), .A1 (n_3443), .A2 (n_2146));
NAND2_X1 i_1110 (.ZN (n_2053), .A1 (inputB[31]), .A2 (inputA[8]));
NOR2_X1 i_1109 (.ZN (n_2052), .A1 (n_3444), .A2 (n_2144));
NAND2_X1 i_1108 (.ZN (n_2051), .A1 (n_2053), .A2 (n_2052));
OAI21_X1 i_1107 (.ZN (n_2050), .A (n_2051), .B1 (n_2053), .B2 (n_2052));
XNOR2_X1 i_1106 (.ZN (n_2049), .A (n_2054), .B (n_2050));
OAI21_X1 i_1105 (.ZN (n_2048), .A (n_2054), .B1 (n_2053), .B2 (n_2052));
NAND2_X1 i_1104 (.ZN (n_2047), .A1 (n_2051), .A2 (n_2048));
NAND2_X1 i_1103 (.ZN (n_2046), .A1 (inputB[10]), .A2 (inputA[30]));
NOR3_X1 i_1102 (.ZN (n_2045), .A1 (n_3420), .A2 (n_3405), .A3 (n_2046));
INV_X1 i_1101 (.ZN (n_2044), .A (n_2045));
AOI22_X1 i_1100 (.ZN (n_2043), .A1 (inputB[10]), .A2 (inputA[29]), .B1 (inputB[9]), .B2 (inputA[30]));
NOR2_X1 i_1099 (.ZN (n_2042), .A1 (n_2045), .A2 (n_2043));
NOR2_X1 i_1098 (.ZN (n_2041), .A1 (n_3419), .A2 (n_3410));
XNOR2_X1 i_1097 (.ZN (n_2040), .A (n_2042), .B (n_2041));
NOR2_X1 i_1096 (.ZN (n_2039), .A1 (n_3443), .A2 (n_2148));
NAND2_X1 i_1095 (.ZN (n_2038), .A1 (inputB[31]), .A2 (inputA[9]));
NOR2_X1 i_1094 (.ZN (n_2037), .A1 (n_3444), .A2 (n_2146));
NAND2_X1 i_1093 (.ZN (n_2036), .A1 (n_2038), .A2 (n_2037));
OAI21_X1 i_1092 (.ZN (n_2035), .A (n_2036), .B1 (n_2038), .B2 (n_2037));
XNOR2_X1 i_1091 (.ZN (n_2034), .A (n_2039), .B (n_2035));
OAI21_X1 i_1090 (.ZN (n_2033), .A (n_2039), .B1 (n_2038), .B2 (n_2037));
NAND2_X1 i_1089 (.ZN (n_2032), .A1 (n_2036), .A2 (n_2033));
NOR2_X1 i_1088 (.ZN (n_2031), .A1 (n_3420), .A2 (n_3410));
NOR2_X1 i_1087 (.ZN (n_2030), .A1 (n_2046), .A2 (n_2031));
AOI21_X1 i_1086 (.ZN (n_2029), .A (n_2030), .B1 (n_2046), .B2 (n_2031));
OAI21_X1 i_1085 (.ZN (n_2028), .A (n_2044), .B1 (n_2043), .B2 (n_2041));
XOR2_X1 i_1084 (.Z (n_2027), .A (n_2029), .B (n_2028));
NOR2_X1 i_1083 (.ZN (n_2026), .A1 (n_2030), .A2 (n_2028));
AOI21_X1 i_1082 (.ZN (n_2025), .A (n_2026), .B1 (n_2046), .B2 (n_2031));
NOR2_X1 i_1081 (.ZN (n_2024), .A1 (n_3443), .A2 (n_2149));
NAND2_X1 i_1080 (.ZN (n_2023), .A1 (inputB[31]), .A2 (inputA[10]));
NOR2_X1 i_1079 (.ZN (n_2022), .A1 (n_3444), .A2 (n_2148));
NAND2_X1 i_1078 (.ZN (n_2021), .A1 (n_2023), .A2 (n_2022));
OAI21_X1 i_1077 (.ZN (n_2020), .A (n_2021), .B1 (n_2023), .B2 (n_2022));
XNOR2_X1 i_1076 (.ZN (n_2019), .A (n_2024), .B (n_2020));
OAI21_X1 i_1075 (.ZN (n_2018), .A (n_2024), .B1 (n_2023), .B2 (n_2022));
NAND2_X1 i_1074 (.ZN (n_2017), .A1 (n_2021), .A2 (n_2018));
NAND2_X1 i_1073 (.ZN (n_2016), .A1 (inputB[10]), .A2 (inputA[31]));
AND2_X1 i_1072 (.ZN (n_2015), .A1 (n_1327), .A2 (n_2016));
NOR2_X1 i_1071 (.ZN (n_2014), .A1 (n_1327), .A2 (n_2016));
NOR2_X1 i_1070 (.ZN (n_2013), .A1 (n_2015), .A2 (n_2014));
XOR2_X1 i_1069 (.Z (n_2012), .A (n_1329), .B (n_2013));
NOR2_X1 i_1068 (.ZN (n_2011), .A1 (n_1329), .A2 (n_2015));
NOR2_X1 i_1067 (.ZN (n_2010), .A1 (n_2014), .A2 (n_2011));
NOR2_X1 i_1066 (.ZN (n_2009), .A1 (n_3443), .A2 (n_2150));
NAND2_X1 i_1065 (.ZN (n_2008), .A1 (inputB[31]), .A2 (inputA[11]));
NOR2_X1 i_1064 (.ZN (n_2007), .A1 (n_3444), .A2 (n_2149));
NAND2_X1 i_1063 (.ZN (n_2006), .A1 (n_2008), .A2 (n_2007));
OAI21_X1 i_1062 (.ZN (n_2005), .A (n_2006), .B1 (n_2008), .B2 (n_2007));
XNOR2_X1 i_1061 (.ZN (n_2004), .A (n_2009), .B (n_2005));
OAI21_X1 i_1060 (.ZN (n_2003), .A (n_2009), .B1 (n_2008), .B2 (n_2007));
NAND2_X1 i_1059 (.ZN (n_2002), .A1 (n_2006), .A2 (n_2003));
NAND2_X1 i_1058 (.ZN (n_2001), .A1 (inputB[13]), .A2 (inputA[30]));
NOR3_X1 i_1057 (.ZN (n_2000), .A1 (n_3426), .A2 (n_3405), .A3 (n_2001));
AOI22_X1 i_1056 (.ZN (n_1999), .A1 (inputB[13]), .A2 (inputA[29]), .B1 (inputB[12]), .B2 (inputA[30]));
NOR2_X1 i_1055 (.ZN (n_1998), .A1 (n_2000), .A2 (n_1999));
NOR2_X1 i_1054 (.ZN (n_1997), .A1 (n_3422), .A2 (n_3410));
NOR2_X1 i_1053 (.ZN (n_1996), .A1 (n_1999), .A2 (n_1997));
XNOR2_X1 i_1052 (.ZN (n_1995), .A (n_1998), .B (n_1997));
NOR2_X1 i_1051 (.ZN (n_1994), .A1 (n_3443), .A2 (n_2151));
NAND2_X1 i_1050 (.ZN (n_1993), .A1 (inputB[31]), .A2 (inputA[12]));
NOR2_X1 i_1049 (.ZN (n_1992), .A1 (n_3444), .A2 (n_2150));
NAND2_X1 i_1048 (.ZN (n_1991), .A1 (n_1993), .A2 (n_1992));
OAI21_X1 i_1047 (.ZN (n_1990), .A (n_1991), .B1 (n_1993), .B2 (n_1992));
XNOR2_X1 i_1046 (.ZN (n_1989), .A (n_1994), .B (n_1990));
OAI21_X1 i_1045 (.ZN (n_1988), .A (n_1994), .B1 (n_1993), .B2 (n_1992));
NAND2_X1 i_1044 (.ZN (n_1987), .A1 (n_1991), .A2 (n_1988));
NOR2_X1 i_1043 (.ZN (n_1986), .A1 (n_3426), .A2 (n_3410));
NAND2_X1 i_1042 (.ZN (n_1985), .A1 (n_2001), .A2 (n_1986));
INV_X1 i_1041 (.ZN (n_1984), .A (n_1985));
OAI21_X1 i_1040 (.ZN (n_1983), .A (n_1985), .B1 (n_2001), .B2 (n_1986));
NOR2_X1 i_1039 (.ZN (n_1982), .A1 (n_2000), .A2 (n_1996));
XOR2_X1 i_1038 (.Z (n_1981), .A (n_1983), .B (n_1982));
OAI22_X1 i_1037 (.ZN (n_1980), .A1 (n_2001), .A2 (n_1986), .B1 (n_1984), .B2 (n_1982));
NOR2_X1 i_1036 (.ZN (n_1979), .A1 (n_3443), .A2 (n_2152));
NAND2_X1 i_1035 (.ZN (n_1978), .A1 (inputB[31]), .A2 (inputA[13]));
NOR2_X1 i_1034 (.ZN (n_1977), .A1 (n_3444), .A2 (n_2151));
NAND2_X1 i_1033 (.ZN (n_1976), .A1 (n_1978), .A2 (n_1977));
OAI21_X1 i_1032 (.ZN (n_1975), .A (n_1976), .B1 (n_1978), .B2 (n_1977));
XNOR2_X1 i_1031 (.ZN (n_1974), .A (n_1979), .B (n_1975));
OAI21_X1 i_1030 (.ZN (n_1973), .A (n_1979), .B1 (n_1978), .B2 (n_1977));
NAND2_X1 i_1029 (.ZN (n_1972), .A1 (n_1976), .A2 (n_1973));
NAND2_X1 i_1028 (.ZN (n_1971), .A1 (inputB[13]), .A2 (inputA[31]));
AND2_X1 i_1027 (.ZN (n_1970), .A1 (n_1439), .A2 (n_1971));
NOR2_X1 i_1026 (.ZN (n_1969), .A1 (n_1439), .A2 (n_1971));
NOR2_X1 i_1025 (.ZN (n_1968), .A1 (n_1970), .A2 (n_1969));
XOR2_X1 i_1024 (.Z (n_1967), .A (n_1441), .B (n_1968));
NOR2_X1 i_1023 (.ZN (n_1966), .A1 (n_1441), .A2 (n_1970));
NOR2_X1 i_1022 (.ZN (n_1965), .A1 (n_1969), .A2 (n_1966));
NOR2_X1 i_1021 (.ZN (n_1964), .A1 (n_3443), .A2 (n_2154));
NAND2_X1 i_1020 (.ZN (n_1963), .A1 (inputB[31]), .A2 (inputA[14]));
NOR2_X1 i_1019 (.ZN (n_1962), .A1 (n_3444), .A2 (n_2152));
NAND2_X1 i_1018 (.ZN (n_1961), .A1 (n_1963), .A2 (n_1962));
OAI21_X1 i_1017 (.ZN (n_1960), .A (n_1961), .B1 (n_1963), .B2 (n_1962));
XNOR2_X1 i_1016 (.ZN (n_1959), .A (n_1964), .B (n_1960));
OAI21_X1 i_1015 (.ZN (n_1958), .A (n_1964), .B1 (n_1963), .B2 (n_1962));
NAND2_X1 i_1014 (.ZN (n_1957), .A1 (n_1961), .A2 (n_1958));
NAND2_X1 i_1013 (.ZN (n_1956), .A1 (inputB[16]), .A2 (inputA[30]));
NOR3_X1 i_1012 (.ZN (n_1955), .A1 (n_3429), .A2 (n_3405), .A3 (n_1956));
INV_X1 i_1011 (.ZN (n_1954), .A (n_1955));
AOI22_X1 i_1010 (.ZN (n_1953), .A1 (inputB[16]), .A2 (inputA[29]), .B1 (inputB[15]), .B2 (inputA[30]));
NOR2_X1 i_1009 (.ZN (n_1952), .A1 (n_1955), .A2 (n_1953));
NOR2_X1 i_1008 (.ZN (n_1951), .A1 (n_3428), .A2 (n_3410));
XNOR2_X1 i_1007 (.ZN (n_1950), .A (n_1952), .B (n_1951));
NOR2_X1 i_1006 (.ZN (n_1949), .A1 (n_3443), .A2 (n_2155));
NAND2_X1 i_1005 (.ZN (n_1948), .A1 (inputB[31]), .A2 (inputA[15]));
NOR2_X1 i_1004 (.ZN (n_1947), .A1 (n_3444), .A2 (n_2154));
NAND2_X1 i_1003 (.ZN (n_1946), .A1 (n_1948), .A2 (n_1947));
OAI21_X1 i_1002 (.ZN (n_1945), .A (n_1946), .B1 (n_1948), .B2 (n_1947));
XNOR2_X1 i_1001 (.ZN (n_1944), .A (n_1949), .B (n_1945));
OAI21_X1 i_1000 (.ZN (n_1943), .A (n_1949), .B1 (n_1948), .B2 (n_1947));
NAND2_X1 i_999 (.ZN (n_1942), .A1 (n_1946), .A2 (n_1943));
NOR2_X1 i_998 (.ZN (n_1941), .A1 (n_3429), .A2 (n_3410));
NOR2_X1 i_997 (.ZN (n_1940), .A1 (n_1956), .A2 (n_1941));
AOI21_X1 i_996 (.ZN (n_1939), .A (n_1940), .B1 (n_1956), .B2 (n_1941));
OAI21_X1 i_995 (.ZN (n_1938), .A (n_1954), .B1 (n_1953), .B2 (n_1951));
XOR2_X1 i_994 (.Z (n_1937), .A (n_1939), .B (n_1938));
NOR2_X1 i_993 (.ZN (n_1936), .A1 (n_1940), .A2 (n_1938));
AOI21_X1 i_992 (.ZN (n_1935), .A (n_1936), .B1 (n_1956), .B2 (n_1941));
NOR2_X1 i_991 (.ZN (n_1934), .A1 (n_3443), .A2 (n_2156));
NAND2_X1 i_990 (.ZN (n_1933), .A1 (inputB[31]), .A2 (inputA[16]));
NOR2_X1 i_989 (.ZN (n_1932), .A1 (n_3444), .A2 (n_2155));
NAND2_X1 i_988 (.ZN (n_1931), .A1 (n_1933), .A2 (n_1932));
OAI21_X1 i_987 (.ZN (n_1930), .A (n_1931), .B1 (n_1933), .B2 (n_1932));
XNOR2_X1 i_986 (.ZN (n_1929), .A (n_1934), .B (n_1930));
OAI21_X1 i_985 (.ZN (n_1928), .A (n_1934), .B1 (n_1933), .B2 (n_1932));
NAND2_X1 i_984 (.ZN (n_1927), .A1 (n_1931), .A2 (n_1928));
NAND2_X1 i_983 (.ZN (n_1926), .A1 (inputB[16]), .A2 (inputA[31]));
AND2_X1 i_982 (.ZN (n_1925), .A1 (n_1533), .A2 (n_1926));
NOR2_X1 i_981 (.ZN (n_1924), .A1 (n_1533), .A2 (n_1926));
NOR2_X1 i_980 (.ZN (n_1923), .A1 (n_1925), .A2 (n_1924));
XOR2_X1 i_979 (.Z (n_1922), .A (n_1535), .B (n_1923));
NOR2_X1 i_978 (.ZN (n_1921), .A1 (n_1535), .A2 (n_1925));
NOR2_X1 i_977 (.ZN (n_1920), .A1 (n_1924), .A2 (n_1921));
NOR2_X1 i_976 (.ZN (n_1919), .A1 (n_3443), .A2 (n_2158));
NAND2_X1 i_975 (.ZN (n_1918), .A1 (inputB[31]), .A2 (inputA[17]));
NOR2_X1 i_974 (.ZN (n_1917), .A1 (n_3444), .A2 (n_2156));
NAND2_X1 i_973 (.ZN (n_1916), .A1 (n_1918), .A2 (n_1917));
OAI21_X1 i_972 (.ZN (n_1915), .A (n_1916), .B1 (n_1918), .B2 (n_1917));
XNOR2_X1 i_971 (.ZN (n_1914), .A (n_1919), .B (n_1915));
OAI21_X1 i_970 (.ZN (n_1913), .A (n_1919), .B1 (n_1918), .B2 (n_1917));
NAND2_X1 i_969 (.ZN (n_1912), .A1 (n_1916), .A2 (n_1913));
NAND2_X1 i_968 (.ZN (n_1911), .A1 (inputB[19]), .A2 (inputA[30]));
NOR3_X1 i_967 (.ZN (n_1910), .A1 (n_3432), .A2 (n_3405), .A3 (n_1911));
INV_X1 i_966 (.ZN (n_1909), .A (n_1910));
AOI22_X1 i_965 (.ZN (n_1908), .A1 (inputB[19]), .A2 (inputA[29]), .B1 (inputB[18]), .B2 (inputA[30]));
NOR2_X1 i_964 (.ZN (n_1907), .A1 (n_1910), .A2 (n_1908));
NOR2_X1 i_963 (.ZN (n_1906), .A1 (n_3431), .A2 (n_3410));
XNOR2_X1 i_962 (.ZN (n_1905), .A (n_1907), .B (n_1906));
NOR2_X1 i_961 (.ZN (n_1904), .A1 (n_3443), .A2 (n_2162));
NAND2_X1 i_960 (.ZN (n_1903), .A1 (inputB[31]), .A2 (inputA[18]));
NOR2_X1 i_959 (.ZN (n_1902), .A1 (n_3444), .A2 (n_2158));
NAND2_X1 i_958 (.ZN (n_1901), .A1 (n_1903), .A2 (n_1902));
OAI21_X1 i_957 (.ZN (n_1900), .A (n_1901), .B1 (n_1903), .B2 (n_1902));
XNOR2_X1 i_956 (.ZN (n_1899), .A (n_1904), .B (n_1900));
OAI21_X1 i_955 (.ZN (n_1898), .A (n_1904), .B1 (n_1903), .B2 (n_1902));
NAND2_X1 i_954 (.ZN (n_1897), .A1 (n_1901), .A2 (n_1898));
NOR2_X1 i_953 (.ZN (n_1896), .A1 (n_3432), .A2 (n_3410));
NOR2_X1 i_952 (.ZN (n_1895), .A1 (n_1911), .A2 (n_1896));
AOI21_X1 i_951 (.ZN (n_1894), .A (n_1895), .B1 (n_1911), .B2 (n_1896));
OAI21_X1 i_950 (.ZN (n_1893), .A (n_1909), .B1 (n_1908), .B2 (n_1906));
XOR2_X1 i_949 (.Z (n_1892), .A (n_1894), .B (n_1893));
NOR2_X1 i_948 (.ZN (n_1891), .A1 (n_1895), .A2 (n_1893));
AOI21_X1 i_947 (.ZN (n_1890), .A (n_1891), .B1 (n_1911), .B2 (n_1896));
NOR2_X1 i_946 (.ZN (n_1889), .A1 (n_3443), .A2 (n_2163));
NAND2_X1 i_945 (.ZN (n_1888), .A1 (inputB[31]), .A2 (inputA[19]));
NOR2_X1 i_944 (.ZN (n_1887), .A1 (n_3444), .A2 (n_2162));
NAND2_X1 i_943 (.ZN (n_1886), .A1 (n_1888), .A2 (n_1887));
OAI21_X1 i_942 (.ZN (n_1885), .A (n_1886), .B1 (n_1888), .B2 (n_1887));
XNOR2_X1 i_941 (.ZN (n_1884), .A (n_1889), .B (n_1885));
OAI21_X1 i_940 (.ZN (n_1883), .A (n_1889), .B1 (n_1888), .B2 (n_1887));
NAND2_X1 i_939 (.ZN (n_1882), .A1 (n_1886), .A2 (n_1883));
NAND2_X1 i_938 (.ZN (n_1881), .A1 (inputB[19]), .A2 (inputA[31]));
AND2_X1 i_937 (.ZN (n_1880), .A1 (n_1609), .A2 (n_1881));
NOR2_X1 i_936 (.ZN (n_1879), .A1 (n_1609), .A2 (n_1881));
NOR2_X1 i_935 (.ZN (n_1878), .A1 (n_1880), .A2 (n_1879));
XOR2_X1 i_934 (.Z (n_1877), .A (n_1611), .B (n_1878));
NOR2_X1 i_933 (.ZN (n_1876), .A1 (n_1611), .A2 (n_1880));
NOR2_X1 i_932 (.ZN (n_1875), .A1 (n_1879), .A2 (n_1876));
NOR2_X1 i_931 (.ZN (n_1874), .A1 (n_3443), .A2 (n_2164));
NAND2_X1 i_930 (.ZN (n_1873), .A1 (inputB[31]), .A2 (inputA[20]));
NOR2_X1 i_929 (.ZN (n_1872), .A1 (n_3444), .A2 (n_2163));
NAND2_X1 i_928 (.ZN (n_1871), .A1 (n_1873), .A2 (n_1872));
OAI21_X1 i_927 (.ZN (n_1870), .A (n_1871), .B1 (n_1873), .B2 (n_1872));
XNOR2_X1 i_926 (.ZN (n_1869), .A (n_1874), .B (n_1870));
OAI21_X1 i_925 (.ZN (n_1868), .A (n_1874), .B1 (n_1873), .B2 (n_1872));
NAND2_X1 i_924 (.ZN (n_1867), .A1 (n_1871), .A2 (n_1868));
NAND2_X1 i_923 (.ZN (n_1866), .A1 (inputB[22]), .A2 (inputA[30]));
NOR3_X1 i_922 (.ZN (n_1865), .A1 (n_3435), .A2 (n_3405), .A3 (n_1866));
AOI22_X1 i_921 (.ZN (n_1864), .A1 (inputB[22]), .A2 (inputA[29]), .B1 (inputB[21]), .B2 (inputA[30]));
NOR2_X1 i_920 (.ZN (n_1863), .A1 (n_1865), .A2 (n_1864));
NOR2_X1 i_919 (.ZN (n_1862), .A1 (n_3434), .A2 (n_3410));
NOR2_X1 i_918 (.ZN (n_1861), .A1 (n_1864), .A2 (n_1862));
XNOR2_X1 i_917 (.ZN (n_1860), .A (n_1863), .B (n_1862));
NOR2_X1 i_916 (.ZN (n_1859), .A1 (n_3443), .A2 (n_2166));
NAND2_X1 i_915 (.ZN (n_1858), .A1 (inputB[31]), .A2 (inputA[21]));
NOR2_X1 i_914 (.ZN (n_1857), .A1 (n_3444), .A2 (n_2164));
NAND2_X1 i_913 (.ZN (n_1856), .A1 (n_1858), .A2 (n_1857));
OAI21_X1 i_912 (.ZN (n_1855), .A (n_1856), .B1 (n_1858), .B2 (n_1857));
XNOR2_X1 i_911 (.ZN (n_1854), .A (n_1859), .B (n_1855));
OAI21_X1 i_910 (.ZN (n_1853), .A (n_1859), .B1 (n_1858), .B2 (n_1857));
NAND2_X1 i_909 (.ZN (n_1852), .A1 (n_1856), .A2 (n_1853));
NOR2_X1 i_908 (.ZN (n_1851), .A1 (n_3435), .A2 (n_3410));
NAND2_X1 i_907 (.ZN (n_1850), .A1 (n_1866), .A2 (n_1851));
INV_X1 i_906 (.ZN (n_1849), .A (n_1850));
OAI21_X1 i_905 (.ZN (n_1848), .A (n_1850), .B1 (n_1866), .B2 (n_1851));
NOR2_X1 i_904 (.ZN (n_1847), .A1 (n_1865), .A2 (n_1861));
XOR2_X1 i_903 (.Z (n_1846), .A (n_1848), .B (n_1847));
OAI22_X1 i_902 (.ZN (n_1845), .A1 (n_1866), .A2 (n_1851), .B1 (n_1849), .B2 (n_1847));
NOR2_X1 i_901 (.ZN (n_1844), .A1 (n_3443), .A2 (n_2169));
NAND2_X1 i_900 (.ZN (n_1843), .A1 (inputB[31]), .A2 (inputA[22]));
NOR2_X1 i_899 (.ZN (n_1842), .A1 (n_3444), .A2 (n_2166));
NAND2_X1 i_898 (.ZN (n_1841), .A1 (n_1843), .A2 (n_1842));
OAI21_X1 i_897 (.ZN (n_1840), .A (n_1841), .B1 (n_1843), .B2 (n_1842));
XNOR2_X1 i_896 (.ZN (n_1839), .A (n_1844), .B (n_1840));
OAI21_X1 i_895 (.ZN (n_1838), .A (n_1844), .B1 (n_1843), .B2 (n_1842));
NAND2_X1 i_894 (.ZN (n_1837), .A1 (n_1841), .A2 (n_1838));
NAND2_X1 i_893 (.ZN (n_1836), .A1 (inputB[22]), .A2 (inputA[31]));
AND2_X1 i_892 (.ZN (n_1835), .A1 (n_1667), .A2 (n_1836));
NOR2_X1 i_891 (.ZN (n_1834), .A1 (n_1667), .A2 (n_1836));
NOR2_X1 i_890 (.ZN (n_1833), .A1 (n_1835), .A2 (n_1834));
XOR2_X1 i_889 (.Z (n_1832), .A (n_1669), .B (n_1833));
NOR2_X1 i_888 (.ZN (n_1831), .A1 (n_1669), .A2 (n_1835));
NOR2_X1 i_887 (.ZN (n_1830), .A1 (n_1834), .A2 (n_1831));
NOR2_X1 i_886 (.ZN (n_1829), .A1 (n_3443), .A2 (n_2170));
NAND2_X1 i_885 (.ZN (n_1828), .A1 (inputB[31]), .A2 (inputA[23]));
NOR2_X1 i_884 (.ZN (n_1827), .A1 (n_3444), .A2 (n_2169));
NAND2_X1 i_883 (.ZN (n_1826), .A1 (n_1828), .A2 (n_1827));
OAI21_X1 i_882 (.ZN (n_1825), .A (n_1826), .B1 (n_1828), .B2 (n_1827));
XNOR2_X1 i_881 (.ZN (n_1824), .A (n_1829), .B (n_1825));
OAI21_X1 i_880 (.ZN (n_1823), .A (n_1829), .B1 (n_1828), .B2 (n_1827));
NAND2_X1 i_879 (.ZN (n_1822), .A1 (n_1826), .A2 (n_1823));
NAND2_X1 i_878 (.ZN (n_1821), .A1 (inputB[25]), .A2 (inputA[30]));
NOR3_X1 i_877 (.ZN (n_1820), .A1 (n_3438), .A2 (n_3405), .A3 (n_1821));
INV_X1 i_876 (.ZN (n_1819), .A (n_1820));
AOI22_X1 i_875 (.ZN (n_1818), .A1 (inputB[25]), .A2 (inputA[29]), .B1 (inputB[24]), .B2 (inputA[30]));
NOR2_X1 i_874 (.ZN (n_1817), .A1 (n_1820), .A2 (n_1818));
NOR2_X1 i_873 (.ZN (n_1816), .A1 (n_3437), .A2 (n_3410));
XNOR2_X1 i_872 (.ZN (n_1815), .A (n_1817), .B (n_1816));
NOR2_X1 i_871 (.ZN (n_1814), .A1 (n_3443), .A2 (n_2171));
NAND2_X1 i_870 (.ZN (n_1813), .A1 (inputB[31]), .A2 (inputA[24]));
NOR2_X1 i_869 (.ZN (n_1812), .A1 (n_3444), .A2 (n_2170));
NAND2_X1 i_868 (.ZN (n_1811), .A1 (n_1813), .A2 (n_1812));
INV_X1 i_867 (.ZN (n_1810), .A (n_1811));
OAI21_X1 i_866 (.ZN (n_1809), .A (n_1811), .B1 (n_1813), .B2 (n_1812));
XNOR2_X1 i_865 (.ZN (n_1808), .A (n_1814), .B (n_1809));
NOR2_X1 i_864 (.ZN (n_1807), .A1 (n_3438), .A2 (n_3410));
NOR2_X1 i_863 (.ZN (n_1806), .A1 (n_1821), .A2 (n_1807));
AOI21_X1 i_862 (.ZN (n_1805), .A (n_1806), .B1 (n_1821), .B2 (n_1807));
OAI21_X1 i_861 (.ZN (n_1804), .A (n_1819), .B1 (n_1818), .B2 (n_1816));
XOR2_X1 i_860 (.Z (n_1803), .A (n_1805), .B (n_1804));
NOR2_X1 i_859 (.ZN (n_1802), .A1 (n_1806), .A2 (n_1804));
AOI21_X1 i_858 (.ZN (n_1801), .A (n_1802), .B1 (n_1821), .B2 (n_1807));
NOR2_X1 i_857 (.ZN (n_1800), .A1 (n_3443), .A2 (n_2172));
NAND2_X1 i_856 (.ZN (n_1799), .A1 (inputB[31]), .A2 (inputA[25]));
NOR2_X1 i_855 (.ZN (n_1798), .A1 (n_3444), .A2 (n_2171));
NAND2_X1 i_854 (.ZN (n_1797), .A1 (n_1799), .A2 (n_1798));
OAI21_X1 i_853 (.ZN (n_1796), .A (n_1797), .B1 (n_1799), .B2 (n_1798));
XNOR2_X1 i_852 (.ZN (n_1795), .A (n_1800), .B (n_1796));
OAI21_X1 i_851 (.ZN (n_1794), .A (n_1800), .B1 (n_1799), .B2 (n_1798));
NAND2_X1 i_850 (.ZN (n_1793), .A1 (n_1797), .A2 (n_1794));
NAND2_X1 i_849 (.ZN (n_1792), .A1 (inputB[25]), .A2 (inputA[31]));
NAND2_X1 i_848 (.ZN (n_1791), .A1 (n_1709), .A2 (n_1792));
NOR2_X1 i_847 (.ZN (n_1790), .A1 (n_1709), .A2 (n_1792));
AOI21_X1 i_846 (.ZN (n_1789), .A (n_1790), .B1 (n_1709), .B2 (n_1792));
OAI22_X1 i_845 (.ZN (n_1788), .A1 (n_1813), .A2 (n_1812), .B1 (n_1814), .B2 (n_1810));
XNOR2_X1 i_844 (.ZN (n_1787), .A (n_1789), .B (n_1788));
OAI21_X1 i_843 (.ZN (n_1786), .A (n_1791), .B1 (n_1790), .B2 (n_1788));
NOR2_X1 i_842 (.ZN (n_1785), .A1 (n_3443), .A2 (n_3404));
NAND2_X1 i_841 (.ZN (n_1784), .A1 (inputB[31]), .A2 (inputA[26]));
NOR2_X1 i_840 (.ZN (n_1783), .A1 (n_3444), .A2 (n_2172));
NAND2_X1 i_839 (.ZN (n_1782), .A1 (n_1784), .A2 (n_1783));
OAI21_X1 i_838 (.ZN (n_1781), .A (n_1782), .B1 (n_1784), .B2 (n_1783));
XNOR2_X1 i_837 (.ZN (n_1780), .A (n_1785), .B (n_1781));
OAI21_X1 i_836 (.ZN (n_1779), .A (n_1785), .B1 (n_1784), .B2 (n_1783));
NAND2_X1 i_835 (.ZN (n_1778), .A1 (n_1782), .A2 (n_1779));
NOR2_X1 i_834 (.ZN (n_1774), .A1 (n_3476), .A2 (n_3475));
XNOR2_X1 i_833 (.ZN (n_1771), .A (n_1774), .B (n_3474));
OAI21_X1 i_832 (.ZN (n_1765), .A (n_3466), .B1 (n_3469), .B2 (n_3468));
XNOR2_X1 i_831 (.ZN (n_1764), .A (n_3467), .B (n_1765));
OAI21_X1 i_830 (.ZN (n_1760), .A (n_3478), .B1 (n_3480), .B2 (n_3479));
XOR2_X1 i_829 (.Z (n_1758), .A (n_1760), .B (n_3472));
OAI21_X1 i_828 (.ZN (n_1753), .A (n_3483), .B1 (n_3485), .B2 (n_3484));
XNOR2_X1 i_827 (.ZN (n_1752), .A (n_3482), .B (n_1753));
AOI21_X1 i_826 (.ZN (n_1745), .A (n_3470), .B1 (n_3481), .B2 (n_3471));
XNOR2_X1 i_825 (.ZN (n_1743), .A (n_1745), .B (n_3464));
FA_X1 i_824 (.CO (n_1737), .S (n_1736), .A (n_1752), .B (n_1743), .CI (n_1733));
FA_X1 i_823 (.CO (n_1735), .S (n_1734), .A (n_1727), .B (n_1729), .CI (n_1732));
FA_X1 i_822 (.CO (n_1733), .S (n_1732), .A (n_1778), .B (n_1758), .CI (n_1764));
FA_X1 i_821 (.CO (n_1731), .S (n_1730), .A (n_1721), .B (n_1723), .CI (n_1728));
FA_X1 i_820 (.CO (n_1729), .S (n_1728), .A (n_1771), .B (n_1780), .CI (n_1726));
FA_X1 i_819 (.CO (n_1727), .S (n_1726), .A (n_1719), .B (n_1793), .CI (n_1786));
FA_X1 i_818 (.CO (n_1725), .S (n_1724), .A (n_1720), .B (n_1715), .CI (n_1722));
FA_X1 i_817 (.CO (n_1723), .S (n_1722), .A (n_1711), .B (n_1787), .CI (n_1713));
FA_X1 i_816 (.CO (n_1721), .S (n_1720), .A (n_1801), .B (n_1718), .CI (n_1795));
FA_X1 i_815 (.CO (n_1719), .S (n_1718), .A (n_2177), .B (n_2206), .CI (n_2236));
FA_X1 i_814 (.CO (n_1717), .S (n_1716), .A (n_1712), .B (n_1714), .CI (n_1705));
FA_X1 i_813 (.CO (n_1715), .S (n_1714), .A (n_1710), .B (n_1701), .CI (n_1703));
FA_X1 i_812 (.CO (n_1713), .S (n_1712), .A (n_1803), .B (n_1708), .CI (n_1808));
FA_X1 i_811 (.CO (n_1711), .S (n_1710), .A (n_1697), .B (n_1822), .CI (n_1699));
FA_X1 i_810 (.CO (n_1709), .S (n_1708), .A (n_2178), .B (n_2207), .CI (n_2237));
FA_X1 i_809 (.CO (n_1707), .S (n_1706), .A (n_1691), .B (n_1693), .CI (n_1704));
FA_X1 i_808 (.CO (n_1705), .S (n_1704), .A (n_1689), .B (n_1700), .CI (n_1702));
FA_X1 i_807 (.CO (n_1703), .S (n_1702), .A (n_1824), .B (n_1687), .CI (n_1698));
FA_X1 i_806 (.CO (n_1701), .S (n_1700), .A (n_1830), .B (n_1815), .CI (n_1696));
FA_X1 i_805 (.CO (n_1699), .S (n_1698), .A (n_1685), .B (n_1683), .CI (n_1837));
FA_X1 i_804 (.CO (n_1697), .S (n_1696), .A (n_2179), .B (n_2208), .CI (n_2238));
FA_X1 i_803 (.CO (n_1695), .S (n_1694), .A (n_1690), .B (n_1679), .CI (n_1692));
FA_X1 i_802 (.CO (n_1693), .S (n_1692), .A (n_1675), .B (n_1688), .CI (n_1677));
FA_X1 i_801 (.CO (n_1691), .S (n_1690), .A (n_1832), .B (n_1673), .CI (n_1686));
FA_X1 i_800 (.CO (n_1689), .S (n_1688), .A (n_1684), .B (n_1682), .CI (n_1839));
FA_X1 i_799 (.CO (n_1687), .S (n_1686), .A (n_1852), .B (n_1671), .CI (n_1845));
FA_X1 i_798 (.CO (n_1685), .S (n_1684), .A (n_2267), .B (n_2296), .CI (n_2326));
FA_X1 i_797 (.CO (n_1683), .S (n_1682), .A (n_2180), .B (n_2209), .CI (n_2239));
FA_X1 i_796 (.CO (n_1681), .S (n_1680), .A (n_1676), .B (n_1663), .CI (n_1678));
FA_X1 i_795 (.CO (n_1679), .S (n_1678), .A (n_1674), .B (n_1672), .CI (n_1661));
FA_X1 i_794 (.CO (n_1677), .S (n_1676), .A (n_1657), .B (n_1655), .CI (n_1659));
FA_X1 i_793 (.CO (n_1675), .S (n_1674), .A (n_1666), .B (n_1854), .CI (n_1670));
FA_X1 i_792 (.CO (n_1673), .S (n_1672), .A (n_1653), .B (n_1846), .CI (n_1668));
FA_X1 i_791 (.CO (n_1671), .S (n_1670), .A (n_1651), .B (n_1649), .CI (n_1867));
FA_X1 i_790 (.CO (n_1669), .S (n_1668), .A (n_2268), .B (n_2297), .CI (n_2327));
FA_X1 i_789 (.CO (n_1667), .S (n_1666), .A (n_2181), .B (n_2210), .CI (n_2240));
FA_X1 i_788 (.CO (n_1665), .S (n_1664), .A (n_1660), .B (n_1645), .CI (n_1662));
FA_X1 i_787 (.CO (n_1663), .S (n_1662), .A (n_1656), .B (n_1658), .CI (n_1643));
FA_X1 i_786 (.CO (n_1661), .S (n_1660), .A (n_1654), .B (n_1641), .CI (n_1639));
FA_X1 i_785 (.CO (n_1659), .S (n_1658), .A (n_1635), .B (n_1652), .CI (n_1637));
FA_X1 i_784 (.CO (n_1657), .S (n_1656), .A (n_1650), .B (n_1648), .CI (n_1869));
FA_X1 i_783 (.CO (n_1655), .S (n_1654), .A (n_1882), .B (n_1875), .CI (n_1860));
FA_X1 i_782 (.CO (n_1653), .S (n_1652), .A (n_1633), .B (n_1631), .CI (n_1629));
FA_X1 i_781 (.CO (n_1651), .S (n_1650), .A (n_2269), .B (n_2298), .CI (n_2328));
FA_X1 i_780 (.CO (n_1649), .S (n_1648), .A (n_2182), .B (n_2211), .CI (n_2241));
FA_X1 i_779 (.CO (n_1647), .S (n_1646), .A (n_1625), .B (n_1642), .CI (n_1644));
FA_X1 i_778 (.CO (n_1645), .S (n_1644), .A (n_1621), .B (n_1640), .CI (n_1623));
FA_X1 i_777 (.CO (n_1643), .S (n_1642), .A (n_1619), .B (n_1638), .CI (n_1636));
FA_X1 i_776 (.CO (n_1641), .S (n_1640), .A (n_1877), .B (n_1617), .CI (n_1615));
FA_X1 i_775 (.CO (n_1639), .S (n_1638), .A (n_1628), .B (n_1884), .CI (n_1634));
FA_X1 i_774 (.CO (n_1637), .S (n_1636), .A (n_1890), .B (n_1632), .CI (n_1630));
FA_X1 i_773 (.CO (n_1635), .S (n_1634), .A (n_1607), .B (n_1897), .CI (n_1613));
FA_X1 i_772 (.CO (n_1633), .S (n_1632), .A (n_2357), .B (n_2386), .CI (n_2416));
FA_X1 i_771 (.CO (n_1631), .S (n_1630), .A (n_2270), .B (n_2299), .CI (n_2329));
FA_X1 i_770 (.CO (n_1629), .S (n_1628), .A (n_2183), .B (n_2212), .CI (n_2242));
FA_X1 i_769 (.CO (n_1627), .S (n_1626), .A (n_1622), .B (n_1603), .CI (n_1624));
FA_X1 i_768 (.CO (n_1625), .S (n_1624), .A (n_1599), .B (n_1620), .CI (n_1601));
FA_X1 i_767 (.CO (n_1623), .S (n_1622), .A (n_1597), .B (n_1616), .CI (n_1618));
FA_X1 i_766 (.CO (n_1621), .S (n_1620), .A (n_1595), .B (n_1593), .CI (n_1614));
FA_X1 i_765 (.CO (n_1619), .S (n_1618), .A (n_1899), .B (n_1591), .CI (n_1612));
FA_X1 i_764 (.CO (n_1617), .S (n_1616), .A (n_1610), .B (n_1608), .CI (n_1606));
FA_X1 i_763 (.CO (n_1615), .S (n_1614), .A (n_1912), .B (n_1589), .CI (n_1892));
FA_X1 i_762 (.CO (n_1613), .S (n_1612), .A (n_1587), .B (n_1585), .CI (n_1583));
FA_X1 i_761 (.CO (n_1611), .S (n_1610), .A (n_2358), .B (n_2387), .CI (n_2417));
FA_X1 i_760 (.CO (n_1609), .S (n_1608), .A (n_2271), .B (n_2300), .CI (n_2330));
FA_X1 i_759 (.CO (n_1607), .S (n_1606), .A (n_2184), .B (n_2213), .CI (n_2243));
FA_X1 i_758 (.CO (n_1605), .S (n_1604), .A (n_1600), .B (n_1579), .CI (n_1602));
FA_X1 i_757 (.CO (n_1603), .S (n_1602), .A (n_1596), .B (n_1598), .CI (n_1577));
FA_X1 i_756 (.CO (n_1601), .S (n_1600), .A (n_1594), .B (n_1592), .CI (n_1575));
FA_X1 i_755 (.CO (n_1599), .S (n_1598), .A (n_1567), .B (n_1573), .CI (n_1571));
FA_X1 i_754 (.CO (n_1597), .S (n_1596), .A (n_1590), .B (n_1588), .CI (n_1569));
FA_X1 i_753 (.CO (n_1595), .S (n_1594), .A (n_1584), .B (n_1582), .CI (n_1914));
FA_X1 i_752 (.CO (n_1593), .S (n_1592), .A (n_1920), .B (n_1905), .CI (n_1586));
FA_X1 i_751 (.CO (n_1591), .S (n_1590), .A (n_1557), .B (n_1927), .CI (n_1565));
FA_X1 i_750 (.CO (n_1589), .S (n_1588), .A (n_1563), .B (n_1561), .CI (n_1559));
FA_X1 i_749 (.CO (n_1587), .S (n_1586), .A (n_2359), .B (n_2388), .CI (n_2418));
FA_X1 i_748 (.CO (n_1585), .S (n_1584), .A (n_2272), .B (n_2301), .CI (n_2331));
FA_X1 i_747 (.CO (n_1583), .S (n_1582), .A (n_2185), .B (n_2214), .CI (n_2244));
FA_X1 i_746 (.CO (n_1581), .S (n_1580), .A (n_1576), .B (n_1553), .CI (n_1578));
FA_X1 i_745 (.CO (n_1579), .S (n_1578), .A (n_1549), .B (n_1574), .CI (n_1551));
FA_X1 i_744 (.CO (n_1577), .S (n_1576), .A (n_1568), .B (n_1570), .CI (n_1572));
FA_X1 i_743 (.CO (n_1575), .S (n_1574), .A (n_1566), .B (n_1545), .CI (n_1547));
FA_X1 i_742 (.CO (n_1573), .S (n_1572), .A (n_1922), .B (n_1543), .CI (n_1541));
FA_X1 i_741 (.CO (n_1571), .S (n_1570), .A (n_1929), .B (n_1539), .CI (n_1564));
FA_X1 i_740 (.CO (n_1569), .S (n_1568), .A (n_1560), .B (n_1558), .CI (n_1556));
FA_X1 i_739 (.CO (n_1567), .S (n_1566), .A (n_1537), .B (n_1935), .CI (n_1562));
FA_X1 i_738 (.CO (n_1565), .S (n_1564), .A (n_1531), .B (n_1529), .CI (n_1942));
FA_X1 i_737 (.CO (n_1563), .S (n_1562), .A (n_2447), .B (n_2476), .CI (n_2506));
FA_X1 i_736 (.CO (n_1561), .S (n_1560), .A (n_2360), .B (n_2389), .CI (n_2419));
FA_X1 i_735 (.CO (n_1559), .S (n_1558), .A (n_2273), .B (n_2302), .CI (n_2332));
FA_X1 i_734 (.CO (n_1557), .S (n_1556), .A (n_2186), .B (n_2215), .CI (n_2245));
FA_X1 i_733 (.CO (n_1555), .S (n_1554), .A (n_1550), .B (n_1525), .CI (n_1552));
FA_X1 i_732 (.CO (n_1553), .S (n_1552), .A (n_1521), .B (n_1548), .CI (n_1523));
FA_X1 i_731 (.CO (n_1551), .S (n_1550), .A (n_1519), .B (n_1546), .CI (n_1544));
FA_X1 i_730 (.CO (n_1549), .S (n_1548), .A (n_1517), .B (n_1542), .CI (n_1540));
FA_X1 i_729 (.CO (n_1547), .S (n_1546), .A (n_1513), .B (n_1511), .CI (n_1515));
FA_X1 i_728 (.CO (n_1545), .S (n_1544), .A (n_1944), .B (n_1538), .CI (n_1536));
FA_X1 i_727 (.CO (n_1543), .S (n_1542), .A (n_1532), .B (n_1530), .CI (n_1528));
FA_X1 i_726 (.CO (n_1541), .S (n_1540), .A (n_1507), .B (n_1937), .CI (n_1534));
FA_X1 i_725 (.CO (n_1539), .S (n_1538), .A (n_1499), .B (n_1957), .CI (n_1509));
FA_X1 i_724 (.CO (n_1537), .S (n_1536), .A (n_1505), .B (n_1503), .CI (n_1501));
FA_X1 i_723 (.CO (n_1535), .S (n_1534), .A (n_2448), .B (n_2477), .CI (n_2507));
FA_X1 i_722 (.CO (n_1533), .S (n_1532), .A (n_2361), .B (n_2390), .CI (n_2420));
FA_X1 i_721 (.CO (n_1531), .S (n_1530), .A (n_2274), .B (n_2303), .CI (n_2333));
FA_X1 i_720 (.CO (n_1529), .S (n_1528), .A (n_2187), .B (n_2216), .CI (n_2246));
FA_X1 i_719 (.CO (n_1527), .S (n_1526), .A (n_1522), .B (n_1495), .CI (n_1524));
FA_X1 i_718 (.CO (n_1525), .S (n_1524), .A (n_1491), .B (n_1520), .CI (n_1493));
FA_X1 i_717 (.CO (n_1523), .S (n_1522), .A (n_1516), .B (n_1489), .CI (n_1518));
FA_X1 i_716 (.CO (n_1521), .S (n_1520), .A (n_1485), .B (n_1514), .CI (n_1512));
FA_X1 i_715 (.CO (n_1519), .S (n_1518), .A (n_1481), .B (n_1510), .CI (n_1487));
FA_X1 i_714 (.CO (n_1517), .S (n_1516), .A (n_1508), .B (n_1506), .CI (n_1483));
FA_X1 i_713 (.CO (n_1515), .S (n_1514), .A (n_1498), .B (n_1959), .CI (n_1479));
FA_X1 i_712 (.CO (n_1513), .S (n_1512), .A (n_1504), .B (n_1502), .CI (n_1500));
FA_X1 i_711 (.CO (n_1511), .S (n_1510), .A (n_1477), .B (n_1965), .CI (n_1950));
FA_X1 i_710 (.CO (n_1509), .S (n_1508), .A (n_1469), .B (n_1467), .CI (n_1972));
FA_X1 i_709 (.CO (n_1507), .S (n_1506), .A (n_1475), .B (n_1473), .CI (n_1471));
FA_X1 i_708 (.CO (n_1505), .S (n_1504), .A (n_2449), .B (n_2478), .CI (n_2508));
FA_X1 i_707 (.CO (n_1503), .S (n_1502), .A (n_2362), .B (n_2391), .CI (n_2421));
FA_X1 i_706 (.CO (n_1501), .S (n_1500), .A (n_2275), .B (n_2304), .CI (n_2334));
FA_X1 i_705 (.CO (n_1499), .S (n_1498), .A (n_2188), .B (n_2217), .CI (n_2247));
FA_X1 i_704 (.CO (n_1497), .S (n_1496), .A (n_1492), .B (n_1463), .CI (n_1494));
FA_X1 i_703 (.CO (n_1495), .S (n_1494), .A (n_1459), .B (n_1490), .CI (n_1461));
FA_X1 i_702 (.CO (n_1493), .S (n_1492), .A (n_1484), .B (n_1457), .CI (n_1488));
FA_X1 i_701 (.CO (n_1491), .S (n_1490), .A (n_1480), .B (n_1455), .CI (n_1486));
FA_X1 i_700 (.CO (n_1489), .S (n_1488), .A (n_1478), .B (n_1453), .CI (n_1482));
FA_X1 i_699 (.CO (n_1487), .S (n_1486), .A (n_1451), .B (n_1449), .CI (n_1447));
FA_X1 i_698 (.CO (n_1485), .S (n_1484), .A (n_1974), .B (n_1476), .CI (n_1967));
FA_X1 i_697 (.CO (n_1483), .S (n_1482), .A (n_1470), .B (n_1468), .CI (n_1466));
FA_X1 i_696 (.CO (n_1481), .S (n_1480), .A (n_1980), .B (n_1474), .CI (n_1472));
FA_X1 i_695 (.CO (n_1479), .S (n_1478), .A (n_1987), .B (n_1445), .CI (n_1443));
FA_X1 i_694 (.CO (n_1477), .S (n_1476), .A (n_1437), .B (n_1435), .CI (n_1433));
FA_X1 i_693 (.CO (n_1475), .S (n_1474), .A (n_2537), .B (n_2566), .CI (n_2596));
FA_X1 i_692 (.CO (n_1473), .S (n_1472), .A (n_2450), .B (n_2479), .CI (n_2509));
FA_X1 i_691 (.CO (n_1471), .S (n_1470), .A (n_2363), .B (n_2392), .CI (n_2422));
FA_X1 i_690 (.CO (n_1469), .S (n_1468), .A (n_2276), .B (n_2305), .CI (n_2335));
FA_X1 i_689 (.CO (n_1467), .S (n_1466), .A (n_2189), .B (n_2218), .CI (n_2248));
FA_X1 i_688 (.CO (n_1465), .S (n_1464), .A (n_1460), .B (n_1429), .CI (n_1462));
FA_X1 i_687 (.CO (n_1463), .S (n_1462), .A (n_1425), .B (n_1458), .CI (n_1427));
FA_X1 i_686 (.CO (n_1461), .S (n_1460), .A (n_1452), .B (n_1423), .CI (n_1456));
FA_X1 i_685 (.CO (n_1459), .S (n_1458), .A (n_1448), .B (n_1421), .CI (n_1454));
FA_X1 i_684 (.CO (n_1457), .S (n_1456), .A (n_1419), .B (n_1417), .CI (n_1450));
FA_X1 i_683 (.CO (n_1455), .S (n_1454), .A (n_1415), .B (n_1413), .CI (n_1446));
FA_X1 i_682 (.CO (n_1453), .S (n_1452), .A (n_1411), .B (n_1444), .CI (n_1442));
FA_X1 i_681 (.CO (n_1451), .S (n_1450), .A (n_1434), .B (n_1432), .CI (n_1989));
FA_X1 i_680 (.CO (n_1449), .S (n_1448), .A (n_1440), .B (n_1438), .CI (n_1436));
FA_X1 i_679 (.CO (n_1447), .S (n_1446), .A (n_1409), .B (n_1407), .CI (n_1981));
FA_X1 i_678 (.CO (n_1445), .S (n_1444), .A (n_1399), .B (n_1397), .CI (n_2002));
FA_X1 i_677 (.CO (n_1443), .S (n_1442), .A (n_1405), .B (n_1403), .CI (n_1401));
FA_X1 i_676 (.CO (n_1441), .S (n_1440), .A (n_2538), .B (n_2567), .CI (n_2597));
FA_X1 i_675 (.CO (n_1439), .S (n_1438), .A (n_2451), .B (n_2480), .CI (n_2510));
FA_X1 i_674 (.CO (n_1437), .S (n_1436), .A (n_2364), .B (n_2393), .CI (n_2423));
FA_X1 i_673 (.CO (n_1435), .S (n_1434), .A (n_2277), .B (n_2306), .CI (n_2336));
FA_X1 i_672 (.CO (n_1433), .S (n_1432), .A (n_2190), .B (n_2219), .CI (n_2249));
FA_X1 i_671 (.CO (n_1431), .S (n_1430), .A (n_1426), .B (n_1393), .CI (n_1428));
FA_X1 i_670 (.CO (n_1429), .S (n_1428), .A (n_1422), .B (n_1424), .CI (n_1391));
FA_X1 i_669 (.CO (n_1427), .S (n_1426), .A (n_1387), .B (n_1420), .CI (n_1389));
FA_X1 i_668 (.CO (n_1425), .S (n_1424), .A (n_1416), .B (n_1385), .CI (n_1418));
FA_X1 i_667 (.CO (n_1423), .S (n_1422), .A (n_1381), .B (n_1414), .CI (n_1412));
FA_X1 i_666 (.CO (n_1421), .S (n_1420), .A (n_1375), .B (n_1410), .CI (n_1383));
FA_X1 i_665 (.CO (n_1419), .S (n_1418), .A (n_1406), .B (n_1379), .CI (n_1377));
FA_X1 i_664 (.CO (n_1417), .S (n_1416), .A (n_2004), .B (n_1373), .CI (n_1408));
FA_X1 i_663 (.CO (n_1415), .S (n_1414), .A (n_1400), .B (n_1398), .CI (n_1396));
FA_X1 i_662 (.CO (n_1413), .S (n_1412), .A (n_1995), .B (n_1404), .CI (n_1402));
FA_X1 i_661 (.CO (n_1411), .S (n_1410), .A (n_2017), .B (n_1371), .CI (n_2010));
FA_X1 i_660 (.CO (n_1409), .S (n_1408), .A (n_1363), .B (n_1361), .CI (n_1359));
FA_X1 i_659 (.CO (n_1407), .S (n_1406), .A (n_1369), .B (n_1367), .CI (n_1365));
FA_X1 i_658 (.CO (n_1405), .S (n_1404), .A (n_2539), .B (n_2568), .CI (n_2598));
FA_X1 i_657 (.CO (n_1403), .S (n_1402), .A (n_2452), .B (n_2481), .CI (n_2511));
FA_X1 i_656 (.CO (n_1401), .S (n_1400), .A (n_2365), .B (n_2394), .CI (n_2424));
FA_X1 i_655 (.CO (n_1399), .S (n_1398), .A (n_2278), .B (n_2307), .CI (n_2337));
FA_X1 i_654 (.CO (n_1397), .S (n_1396), .A (n_2191), .B (n_2220), .CI (n_2250));
FA_X1 i_653 (.CO (n_1395), .S (n_1394), .A (n_1390), .B (n_1355), .CI (n_1392));
FA_X1 i_652 (.CO (n_1393), .S (n_1392), .A (n_1386), .B (n_1353), .CI (n_1388));
FA_X1 i_651 (.CO (n_1391), .S (n_1390), .A (n_1349), .B (n_1384), .CI (n_1351));
FA_X1 i_650 (.CO (n_1389), .S (n_1388), .A (n_1382), .B (n_1380), .CI (n_1347));
FA_X1 i_649 (.CO (n_1387), .S (n_1386), .A (n_1378), .B (n_1376), .CI (n_1345));
FA_X1 i_648 (.CO (n_1385), .S (n_1384), .A (n_1341), .B (n_1374), .CI (n_1343));
FA_X1 i_647 (.CO (n_1383), .S (n_1382), .A (n_2012), .B (n_1339), .CI (n_1337));
FA_X1 i_646 (.CO (n_1381), .S (n_1380), .A (n_1335), .B (n_1372), .CI (n_1370));
FA_X1 i_645 (.CO (n_1379), .S (n_1378), .A (n_1360), .B (n_1358), .CI (n_2019));
FA_X1 i_644 (.CO (n_1377), .S (n_1376), .A (n_1366), .B (n_1364), .CI (n_1362));
FA_X1 i_643 (.CO (n_1375), .S (n_1374), .A (n_1331), .B (n_2025), .CI (n_1368));
FA_X1 i_642 (.CO (n_1373), .S (n_1372), .A (n_1319), .B (n_2032), .CI (n_1333));
FA_X1 i_641 (.CO (n_1371), .S (n_1370), .A (n_1325), .B (n_1323), .CI (n_1321));
FA_X1 i_640 (.CO (n_1369), .S (n_1368), .A (n_2627), .B (n_2656), .CI (n_2686));
FA_X1 i_639 (.CO (n_1367), .S (n_1366), .A (n_2540), .B (n_2569), .CI (n_2599));
FA_X1 i_638 (.CO (n_1365), .S (n_1364), .A (n_2453), .B (n_2482), .CI (n_2512));
FA_X1 i_637 (.CO (n_1363), .S (n_1362), .A (n_2366), .B (n_2395), .CI (n_2425));
FA_X1 i_636 (.CO (n_1361), .S (n_1360), .A (n_2279), .B (n_2308), .CI (n_2338));
FA_X1 i_635 (.CO (n_1359), .S (n_1358), .A (n_2192), .B (n_2221), .CI (n_2251));
FA_X1 i_634 (.CO (n_1357), .S (n_1356), .A (n_1352), .B (n_1315), .CI (n_1354));
FA_X1 i_633 (.CO (n_1355), .S (n_1354), .A (n_1348), .B (n_1350), .CI (n_1313));
FA_X1 i_632 (.CO (n_1353), .S (n_1352), .A (n_1309), .B (n_1346), .CI (n_1311));
FA_X1 i_631 (.CO (n_1351), .S (n_1350), .A (n_1344), .B (n_1342), .CI (n_1307));
FA_X1 i_630 (.CO (n_1349), .S (n_1348), .A (n_1338), .B (n_1336), .CI (n_1305));
FA_X1 i_629 (.CO (n_1347), .S (n_1346), .A (n_1303), .B (n_1301), .CI (n_1340));
FA_X1 i_628 (.CO (n_1345), .S (n_1344), .A (n_1297), .B (n_1295), .CI (n_1334));
FA_X1 i_627 (.CO (n_1343), .S (n_1342), .A (n_1332), .B (n_1330), .CI (n_1299));
FA_X1 i_626 (.CO (n_1341), .S (n_1340), .A (n_1318), .B (n_2034), .CI (n_1293));
FA_X1 i_625 (.CO (n_1339), .S (n_1338), .A (n_1324), .B (n_1322), .CI (n_1320));
FA_X1 i_624 (.CO (n_1337), .S (n_1336), .A (n_2027), .B (n_1328), .CI (n_1326));
FA_X1 i_623 (.CO (n_1335), .S (n_1334), .A (n_2047), .B (n_1291), .CI (n_1289));
FA_X1 i_622 (.CO (n_1333), .S (n_1332), .A (n_1281), .B (n_1279), .CI (n_1277));
FA_X1 i_621 (.CO (n_1331), .S (n_1330), .A (n_1287), .B (n_1285), .CI (n_1283));
FA_X1 i_620 (.CO (n_1329), .S (n_1328), .A (n_2628), .B (n_2657), .CI (n_2687));
FA_X1 i_619 (.CO (n_1327), .S (n_1326), .A (n_2541), .B (n_2570), .CI (n_2600));
FA_X1 i_618 (.CO (n_1325), .S (n_1324), .A (n_2454), .B (n_2483), .CI (n_2513));
FA_X1 i_617 (.CO (n_1323), .S (n_1322), .A (n_2367), .B (n_2396), .CI (n_2426));
FA_X1 i_616 (.CO (n_1321), .S (n_1320), .A (n_2280), .B (n_2309), .CI (n_2339));
FA_X1 i_615 (.CO (n_1319), .S (n_1318), .A (n_2193), .B (n_2222), .CI (n_2252));
FA_X1 i_614 (.CO (n_1317), .S (n_1316), .A (n_1312), .B (n_1273), .CI (n_1314));
FA_X1 i_613 (.CO (n_1315), .S (n_1314), .A (n_1269), .B (n_1310), .CI (n_1271));
FA_X1 i_612 (.CO (n_1313), .S (n_1312), .A (n_1306), .B (n_1267), .CI (n_1308));
FA_X1 i_611 (.CO (n_1311), .S (n_1310), .A (n_1302), .B (n_1265), .CI (n_1304));
FA_X1 i_610 (.CO (n_1309), .S (n_1308), .A (n_1296), .B (n_1300), .CI (n_1263));
FA_X1 i_609 (.CO (n_1307), .S (n_1306), .A (n_1261), .B (n_1259), .CI (n_1298));
FA_X1 i_608 (.CO (n_1305), .S (n_1304), .A (n_1253), .B (n_1257), .CI (n_1294));
FA_X1 i_607 (.CO (n_1303), .S (n_1302), .A (n_1290), .B (n_1288), .CI (n_1255));
FA_X1 i_606 (.CO (n_1301), .S (n_1300), .A (n_2049), .B (n_1251), .CI (n_1292));
FA_X1 i_605 (.CO (n_1299), .S (n_1298), .A (n_1280), .B (n_1278), .CI (n_1276));
FA_X1 i_604 (.CO (n_1297), .S (n_1296), .A (n_1286), .B (n_1284), .CI (n_1282));
FA_X1 i_603 (.CO (n_1295), .S (n_1294), .A (n_1247), .B (n_2055), .CI (n_2040));
FA_X1 i_602 (.CO (n_1293), .S (n_1292), .A (n_1233), .B (n_2062), .CI (n_1249));
FA_X1 i_601 (.CO (n_1291), .S (n_1290), .A (n_1239), .B (n_1237), .CI (n_1235));
FA_X1 i_600 (.CO (n_1289), .S (n_1288), .A (n_1245), .B (n_1243), .CI (n_1241));
FA_X1 i_599 (.CO (n_1287), .S (n_1286), .A (n_2629), .B (n_2658), .CI (n_2688));
FA_X1 i_598 (.CO (n_1285), .S (n_1284), .A (n_2542), .B (n_2571), .CI (n_2601));
FA_X1 i_597 (.CO (n_1283), .S (n_1282), .A (n_2455), .B (n_2484), .CI (n_2514));
FA_X1 i_596 (.CO (n_1281), .S (n_1280), .A (n_2368), .B (n_2397), .CI (n_2427));
FA_X1 i_595 (.CO (n_1279), .S (n_1278), .A (n_2281), .B (n_2310), .CI (n_2340));
FA_X1 i_594 (.CO (n_1277), .S (n_1276), .A (n_2194), .B (n_2223), .CI (n_2253));
FA_X1 i_593 (.CO (n_1275), .S (n_1274), .A (n_1229), .B (n_1270), .CI (n_1272));
FA_X1 i_592 (.CO (n_1273), .S (n_1272), .A (n_1225), .B (n_1268), .CI (n_1227));
FA_X1 i_591 (.CO (n_1271), .S (n_1270), .A (n_1223), .B (n_1264), .CI (n_1266));
FA_X1 i_590 (.CO (n_1269), .S (n_1268), .A (n_1258), .B (n_1221), .CI (n_1262));
FA_X1 i_589 (.CO (n_1267), .S (n_1266), .A (n_1252), .B (n_1219), .CI (n_1260));
FA_X1 i_588 (.CO (n_1265), .S (n_1264), .A (n_1215), .B (n_1256), .CI (n_1254));
FA_X1 i_587 (.CO (n_1263), .S (n_1262), .A (n_1213), .B (n_1250), .CI (n_1217));
FA_X1 i_586 (.CO (n_1261), .S (n_1260), .A (n_1211), .B (n_1209), .CI (n_1207));
FA_X1 i_585 (.CO (n_1259), .S (n_1258), .A (n_1248), .B (n_1246), .CI (n_2057));
FA_X1 i_584 (.CO (n_1257), .S (n_1256), .A (n_1232), .B (n_2064), .CI (n_1205));
FA_X1 i_583 (.CO (n_1255), .S (n_1254), .A (n_1238), .B (n_1236), .CI (n_1234));
FA_X1 i_582 (.CO (n_1253), .S (n_1252), .A (n_1244), .B (n_1242), .CI (n_1240));
FA_X1 i_581 (.CO (n_1251), .S (n_1250), .A (n_1203), .B (n_1201), .CI (n_2070));
FA_X1 i_580 (.CO (n_1249), .S (n_1248), .A (n_1189), .B (n_1187), .CI (n_2077));
FA_X1 i_579 (.CO (n_1247), .S (n_1246), .A (n_1195), .B (n_1193), .CI (n_1191));
FA_X1 i_578 (.CO (n_1245), .S (n_1244), .A (n_2717), .B (n_2746), .CI (n_2776));
FA_X1 i_577 (.CO (n_1243), .S (n_1242), .A (n_2630), .B (n_2659), .CI (n_2689));
FA_X1 i_576 (.CO (n_1241), .S (n_1240), .A (n_2543), .B (n_2572), .CI (n_2602));
FA_X1 i_575 (.CO (n_1239), .S (n_1238), .A (n_2456), .B (n_2485), .CI (n_2515));
FA_X1 i_574 (.CO (n_1237), .S (n_1236), .A (n_2369), .B (n_2398), .CI (n_2428));
FA_X1 i_573 (.CO (n_1235), .S (n_1234), .A (n_2282), .B (n_2311), .CI (n_2341));
FA_X1 i_572 (.CO (n_1233), .S (n_1232), .A (n_2195), .B (n_2224), .CI (n_2254));
FA_X1 i_571 (.CO (n_1231), .S (n_1230), .A (n_1183), .B (n_1226), .CI (n_1228));
FA_X1 i_570 (.CO (n_1229), .S (n_1228), .A (n_1222), .B (n_1224), .CI (n_1181));
FA_X1 i_569 (.CO (n_1227), .S (n_1226), .A (n_1177), .B (n_1220), .CI (n_1179));
FA_X1 i_568 (.CO (n_1225), .S (n_1224), .A (n_1173), .B (n_1175), .CI (n_1218));
FA_X1 i_567 (.CO (n_1223), .S (n_1222), .A (n_1171), .B (n_1216), .CI (n_1214));
FA_X1 i_566 (.CO (n_1221), .S (n_1220), .A (n_1212), .B (n_1210), .CI (n_1208));
FA_X1 i_565 (.CO (n_1219), .S (n_1218), .A (n_1206), .B (n_1169), .CI (n_1167));
FA_X1 i_564 (.CO (n_1217), .S (n_1216), .A (n_1165), .B (n_1163), .CI (n_1161));
FA_X1 i_563 (.CO (n_1215), .S (n_1214), .A (n_1204), .B (n_1202), .CI (n_1200));
FA_X1 i_562 (.CO (n_1213), .S (n_1212), .A (n_1186), .B (n_2079), .CI (n_1159));
FA_X1 i_561 (.CO (n_1211), .S (n_1210), .A (n_1192), .B (n_1190), .CI (n_1188));
FA_X1 i_560 (.CO (n_1209), .S (n_1208), .A (n_1198), .B (n_1196), .CI (n_1194));
FA_X1 i_559 (.CO (n_1207), .S (n_1206), .A (n_1155), .B (n_1153), .CI (n_2071));
FA_X1 i_558 (.CO (n_1205), .S (n_1204), .A (n_1139), .B (n_2092), .CI (n_1157));
FA_X1 i_557 (.CO (n_1203), .S (n_1202), .A (n_1145), .B (n_1143), .CI (n_1141));
FA_X1 i_556 (.CO (n_1201), .S (n_1200), .A (n_1151), .B (n_1149), .CI (n_1147));
FA_X1 i_555 (.CO (n_1199), .S (n_1198), .A (n_2718), .B (n_2747), .CI (n_2777));
FA_X1 i_554 (.CO (n_1197), .S (n_1196), .A (n_2631), .B (n_2660), .CI (n_2690));
FA_X1 i_553 (.CO (n_1195), .S (n_1194), .A (n_2544), .B (n_2573), .CI (n_2603));
FA_X1 i_552 (.CO (n_1193), .S (n_1192), .A (n_2457), .B (n_2486), .CI (n_2516));
FA_X1 i_551 (.CO (n_1191), .S (n_1190), .A (n_2370), .B (n_2399), .CI (n_2429));
FA_X1 i_550 (.CO (n_1189), .S (n_1188), .A (n_2283), .B (n_2312), .CI (n_2342));
FA_X1 i_549 (.CO (n_1187), .S (n_1186), .A (n_2196), .B (n_2225), .CI (n_2255));
FA_X1 i_548 (.CO (n_1185), .S (n_1184), .A (n_1180), .B (n_1135), .CI (n_1182));
FA_X1 i_547 (.CO (n_1183), .S (n_1182), .A (n_1176), .B (n_1178), .CI (n_1133));
FA_X1 i_546 (.CO (n_1181), .S (n_1180), .A (n_1129), .B (n_1174), .CI (n_1131));
FA_X1 i_545 (.CO (n_1179), .S (n_1178), .A (n_1170), .B (n_1127), .CI (n_1172));
FA_X1 i_544 (.CO (n_1177), .S (n_1176), .A (n_1168), .B (n_1166), .CI (n_1125));
FA_X1 i_543 (.CO (n_1175), .S (n_1174), .A (n_1162), .B (n_1160), .CI (n_1123));
FA_X1 i_542 (.CO (n_1173), .S (n_1172), .A (n_1121), .B (n_1119), .CI (n_1164));
FA_X1 i_541 (.CO (n_1171), .S (n_1170), .A (n_1111), .B (n_1117), .CI (n_1158));
FA_X1 i_540 (.CO (n_1169), .S (n_1168), .A (n_1152), .B (n_1115), .CI (n_1113));
FA_X1 i_539 (.CO (n_1167), .S (n_1166), .A (n_1109), .B (n_1156), .CI (n_1154));
FA_X1 i_538 (.CO (n_1165), .S (n_1164), .A (n_1140), .B (n_1138), .CI (n_2094));
FA_X1 i_537 (.CO (n_1163), .S (n_1162), .A (n_1146), .B (n_1144), .CI (n_1142));
FA_X1 i_536 (.CO (n_1161), .S (n_1160), .A (n_2085), .B (n_1150), .CI (n_1148));
FA_X1 i_535 (.CO (n_1159), .S (n_1158), .A (n_1107), .B (n_1105), .CI (n_2100));
FA_X1 i_534 (.CO (n_1157), .S (n_1156), .A (n_1091), .B (n_1089), .CI (n_2107));
FA_X1 i_533 (.CO (n_1155), .S (n_1154), .A (n_1097), .B (n_1095), .CI (n_1093));
FA_X1 i_532 (.CO (n_1153), .S (n_1152), .A (n_1103), .B (n_1101), .CI (n_1099));
FA_X1 i_531 (.CO (n_1151), .S (n_1150), .A (n_2719), .B (n_2748), .CI (n_2778));
FA_X1 i_530 (.CO (n_1149), .S (n_1148), .A (n_2632), .B (n_2661), .CI (n_2691));
FA_X1 i_529 (.CO (n_1147), .S (n_1146), .A (n_2545), .B (n_2574), .CI (n_2604));
FA_X1 i_528 (.CO (n_1145), .S (n_1144), .A (n_2458), .B (n_2487), .CI (n_2517));
FA_X1 i_527 (.CO (n_1143), .S (n_1142), .A (n_2371), .B (n_2400), .CI (n_2430));
FA_X1 i_526 (.CO (n_1141), .S (n_1140), .A (n_2284), .B (n_2313), .CI (n_2343));
FA_X1 i_525 (.CO (n_1139), .S (n_1138), .A (n_2197), .B (n_2226), .CI (n_2256));
FA_X1 i_524 (.CO (n_1137), .S (n_1136), .A (n_1132), .B (n_1085), .CI (n_1134));
FA_X1 i_523 (.CO (n_1135), .S (n_1134), .A (n_1128), .B (n_1083), .CI (n_1130));
FA_X1 i_522 (.CO (n_1133), .S (n_1132), .A (n_1079), .B (n_1126), .CI (n_1081));
FA_X1 i_521 (.CO (n_1131), .S (n_1130), .A (n_1077), .B (n_1124), .CI (n_1122));
FA_X1 i_520 (.CO (n_1129), .S (n_1128), .A (n_1120), .B (n_1118), .CI (n_1075));
FA_X1 i_519 (.CO (n_1127), .S (n_1126), .A (n_1114), .B (n_1112), .CI (n_1073));
FA_X1 i_518 (.CO (n_1125), .S (n_1124), .A (n_1069), .B (n_768), .CI (n_1116));
FA_X1 i_517 (.CO (n_1123), .S (n_1122), .A (n_1110), .B (n_1108), .CI (n_1071));
FA_X1 i_516 (.CO (n_1121), .S (n_1120), .A (n_1065), .B (n_1063), .CI (n_1061));
FA_X1 i_515 (.CO (n_1119), .S (n_1118), .A (n_1106), .B (n_1104), .CI (n_2102));
FA_X1 i_514 (.CO (n_1117), .S (n_1116), .A (n_1088), .B (n_2109), .CI (n_1059));
FA_X1 i_513 (.CO (n_1115), .S (n_1114), .A (n_1094), .B (n_1092), .CI (n_1090));
FA_X1 i_512 (.CO (n_1113), .S (n_1112), .A (n_1100), .B (n_1098), .CI (n_1096));
FA_X1 i_511 (.CO (n_1111), .S (n_1110), .A (n_1053), .B (n_2115), .CI (n_1102));
FA_X1 i_510 (.CO (n_1109), .S (n_1108), .A (n_2122), .B (n_766), .CI (n_1055));
FA_X1 i_509 (.CO (n_1107), .S (n_1106), .A (n_1041), .B (n_1039), .CI (n_1037));
FA_X1 i_508 (.CO (n_1105), .S (n_1104), .A (n_1047), .B (n_1045), .CI (n_1043));
FA_X1 i_507 (.CO (n_1103), .S (n_1102), .A (n_2807), .B (n_2836), .CI (n_2866));
FA_X1 i_506 (.CO (n_1101), .S (n_1100), .A (n_2720), .B (n_2749), .CI (n_2779));
FA_X1 i_505 (.CO (n_1099), .S (n_1098), .A (n_2633), .B (n_2662), .CI (n_2692));
FA_X1 i_504 (.CO (n_1097), .S (n_1096), .A (n_2546), .B (n_2575), .CI (n_2605));
FA_X1 i_503 (.CO (n_1095), .S (n_1094), .A (n_2459), .B (n_2488), .CI (n_2518));
FA_X1 i_502 (.CO (n_1093), .S (n_1092), .A (n_2372), .B (n_2401), .CI (n_2431));
FA_X1 i_501 (.CO (n_1091), .S (n_1090), .A (n_2285), .B (n_2314), .CI (n_2344));
FA_X1 i_500 (.CO (n_1089), .S (n_1088), .A (n_2198), .B (n_2227), .CI (n_2257));
FA_X1 i_499 (.CO (n_1087), .S (n_1086), .A (n_1082), .B (n_1033), .CI (n_1084));
FA_X1 i_498 (.CO (n_1085), .S (n_1084), .A (n_1078), .B (n_1080), .CI (n_1031));
FA_X1 i_497 (.CO (n_1083), .S (n_1082), .A (n_1074), .B (n_1076), .CI (n_1029));
FA_X1 i_496 (.CO (n_1081), .S (n_1080), .A (n_1072), .B (n_1027), .CI (n_1025));
FA_X1 i_495 (.CO (n_1079), .S (n_1078), .A (n_1070), .B (n_1068), .CI (n_1023));
FA_X1 i_494 (.CO (n_1075), .S (n_1074), .A (n_1064), .B (n_1062), .CI (n_1060));
FA_X1 i_493 (.CO (n_1073), .S (n_1072), .A (n_1058), .B (n_1017), .CI (n_1015));
FA_X1 i_492 (.CO (n_1071), .S (n_1070), .A (n_1011), .B (n_1009), .CI (n_1057));
FA_X1 i_491 (.CO (n_1069), .S (n_1068), .A (n_1054), .B (n_1052), .CI (n_1013));
FA_X1 i_490 (.CO (n_1065), .S (n_1064), .A (n_1040), .B (n_1038), .CI (n_1036));
FA_X1 i_489 (.CO (n_1063), .S (n_1062), .A (n_1046), .B (n_1044), .CI (n_1042));
FA_X1 i_488 (.CO (n_1061), .S (n_1060), .A (n_2116), .B (n_1050), .CI (n_1048));
FA_X1 i_487 (.CO (n_1059), .S (n_1058), .A (n_1003), .B (n_1001), .CI (n_999));
FA_X1 i_486 (.CO (n_1055), .S (n_1054), .A (n_991), .B (n_989), .CI (n_987));
FA_X1 i_485 (.CO (n_1053), .S (n_1052), .A (n_997), .B (n_995), .CI (n_993));
FA_X1 i_484 (.CO (n_1051), .S (n_1050), .A (n_2808), .B (n_2837), .CI (n_2867));
FA_X1 i_483 (.CO (n_1049), .S (n_1048), .A (n_2721), .B (n_2750), .CI (n_2780));
FA_X1 i_482 (.CO (n_1047), .S (n_1046), .A (n_2634), .B (n_2663), .CI (n_2693));
FA_X1 i_481 (.CO (n_1045), .S (n_1044), .A (n_2547), .B (n_2576), .CI (n_2606));
FA_X1 i_480 (.CO (n_1043), .S (n_1042), .A (n_2460), .B (n_2489), .CI (n_2519));
FA_X1 i_479 (.CO (n_1041), .S (n_1040), .A (n_2373), .B (n_2402), .CI (n_2432));
FA_X1 i_478 (.CO (n_1039), .S (n_1038), .A (n_2286), .B (n_2315), .CI (n_2345));
FA_X1 i_477 (.CO (n_1037), .S (n_1036), .A (n_2199), .B (n_2228), .CI (n_2258));
FA_X1 i_476 (.CO (n_1035), .S (n_1034), .A (n_1030), .B (n_979), .CI (n_1032));
FA_X1 i_475 (.CO (n_1033), .S (n_1032), .A (n_975), .B (n_1028), .CI (n_977));
FA_X1 i_474 (.CO (n_1031), .S (n_1030), .A (n_1022), .B (n_1026), .CI (n_1024));
FA_X1 i_473 (.CO (n_1029), .S (n_1028), .A (n_943), .B (n_971), .CI (n_973));
FA_X1 i_472 (.CO (n_1027), .S (n_1026), .A (n_1014), .B (n_969), .CI (n_967));
FA_X1 i_471 (.CO (n_1025), .S (n_1024), .A (n_965), .B (n_1067), .CI (n_1016));
FA_X1 i_470 (.CO (n_1023), .S (n_1022), .A (n_1012), .B (n_1010), .CI (n_1008));
FA_X1 i_469 (.CO (n_1017), .S (n_1016), .A (n_998), .B (n_959), .CI (n_957));
FA_X1 i_468 (.CO (n_1015), .S (n_1014), .A (n_951), .B (n_1002), .CI (n_1000));
FA_X1 i_467 (.CO (n_1013), .S (n_1012), .A (n_762), .B (n_764), .CI (n_2139));
FA_X1 i_466 (.CO (n_1011), .S (n_1010), .A (n_990), .B (n_988), .CI (n_986));
FA_X1 i_465 (.CO (n_1009), .S (n_1008), .A (n_996), .B (n_994), .CI (n_992));
FA_X1 i_464 (.CO (n_1003), .S (n_1002), .A (n_931), .B (n_929), .CI (n_927));
FA_X1 i_463 (.CO (n_1001), .S (n_1000), .A (n_960), .B (n_935), .CI (n_933));
FA_X1 i_462 (.CO (n_999), .S (n_998), .A (n_1018), .B (n_952), .CI (n_954));
FA_X1 i_461 (.CO (n_997), .S (n_996), .A (n_2809), .B (n_2838), .CI (n_2868));
FA_X1 i_460 (.CO (n_995), .S (n_994), .A (n_2722), .B (n_2751), .CI (n_2781));
FA_X1 i_459 (.CO (n_993), .S (n_992), .A (n_2635), .B (n_2664), .CI (n_2694));
FA_X1 i_458 (.CO (n_991), .S (n_990), .A (n_2548), .B (n_2577), .CI (n_2607));
FA_X1 i_457 (.CO (n_989), .S (n_988), .A (n_2461), .B (n_2490), .CI (n_2520));
FA_X1 i_456 (.CO (n_987), .S (n_986), .A (n_2374), .B (n_2403), .CI (n_2433));
FA_X1 i_455 (.CO (n_981), .S (n_980), .A (n_976), .B (n_978), .CI (n_923));
FA_X1 i_454 (.CO (n_979), .S (n_978), .A (n_919), .B (n_974), .CI (n_921));
FA_X1 i_453 (.CO (n_977), .S (n_976), .A (n_917), .B (n_970), .CI (n_972));
FA_X1 i_452 (.CO (n_975), .S (n_974), .A (n_966), .B (n_915), .CI (n_968));
FA_X1 i_451 (.CO (n_973), .S (n_972), .A (n_911), .B (n_964), .CI (n_913));
FA_X1 i_450 (.CO (n_971), .S (n_970), .A (n_909), .B (n_830), .CI (n_941));
FA_X1 i_449 (.CO (n_969), .S (n_968), .A (n_956), .B (n_962), .CI (n_1020));
FA_X1 i_448 (.CO (n_967), .S (n_966), .A (n_907), .B (n_905), .CI (n_958));
FA_X1 i_447 (.CO (n_965), .S (n_964), .A (n_897), .B (n_903), .CI (n_950));
FA_X1 i_446 (.CO (n_959), .S (n_958), .A (n_928), .B (n_926), .CI (n_2153));
FA_X1 i_445 (.CO (n_957), .S (n_956), .A (n_934), .B (n_932), .CI (n_930));
FA_X1 i_444 (.CO (n_951), .S (n_950), .A (n_893), .B (n_891), .CI (n_889));
FA_X1 i_443 (.CO (n_935), .S (n_934), .A (n_2521), .B (n_2549), .CI (n_2578));
FA_X1 i_442 (.CO (n_933), .S (n_932), .A (n_2434), .B (n_2462), .CI (n_2491));
FA_X1 i_441 (.CO (n_931), .S (n_930), .A (n_2347), .B (n_2375), .CI (n_2404));
FA_X1 i_440 (.CO (n_929), .S (n_928), .A (n_2260), .B (n_2288), .CI (n_2317));
FA_X1 i_439 (.CO (n_927), .S (n_926), .A (n_2174), .B (n_2201), .CI (n_2230));
HA_X1 i_438 (.CO (n_925), .S (n_924), .A (n_867), .B (n_922));
FA_X1 i_437 (.CO (n_923), .S (n_922), .A (n_865), .B (n_918), .CI (n_920));
FA_X1 i_436 (.CO (n_921), .S (n_920), .A (n_914), .B (n_863), .CI (n_916));
FA_X1 i_435 (.CO (n_919), .S (n_918), .A (n_912), .B (n_910), .CI (n_861));
FA_X1 i_434 (.CO (n_917), .S (n_916), .A (n_857), .B (n_908), .CI (n_859));
FA_X1 i_433 (.CO (n_915), .S (n_914), .A (n_853), .B (n_906), .CI (n_904));
FA_X1 i_432 (.CO (n_913), .S (n_912), .A (n_774), .B (n_896), .CI (n_855));
FA_X1 i_431 (.CO (n_911), .S (n_910), .A (n_849), .B (n_902), .CI (n_772));
FA_X1 i_430 (.CO (n_909), .S (n_908), .A (n_841), .B (n_939), .CI (n_851));
FA_X1 i_429 (.CO (n_907), .S (n_906), .A (n_847), .B (n_845), .CI (n_843));
FA_X1 i_428 (.CO (n_905), .S (n_904), .A (n_892), .B (n_890), .CI (n_888));
FA_X1 i_427 (.CO (n_903), .S (n_902), .A (n_760), .B (n_2167), .CI (n_839));
FA_X1 i_426 (.CO (n_897), .S (n_896), .A (n_2159), .B (n_1007), .CI (n_770));
FA_X1 i_425 (.CO (n_893), .S (n_892), .A (n_817), .B (n_815), .CI (n_813));
FA_X1 i_424 (.CO (n_891), .S (n_890), .A (n_823), .B (n_821), .CI (n_819));
FA_X1 i_423 (.CO (n_889), .S (n_888), .A (n_829), .B (n_827), .CI (n_825));
HA_X1 i_422 (.CO (n_869), .S (n_868), .A (n_809), .B (n_866));
FA_X1 i_421 (.CO (n_867), .S (n_866), .A (n_807), .B (n_862), .CI (n_864));
FA_X1 i_420 (.CO (n_865), .S (n_864), .A (n_860), .B (n_858), .CI (n_805));
FA_X1 i_419 (.CO (n_863), .S (n_862), .A (n_801), .B (n_856), .CI (n_803));
FA_X1 i_418 (.CO (n_861), .S (n_860), .A (n_848), .B (n_799), .CI (n_854));
FA_X1 i_417 (.CO (n_859), .S (n_858), .A (n_797), .B (n_852), .CI (n_850));
FA_X1 i_416 (.CO (n_857), .S (n_856), .A (n_846), .B (n_844), .CI (n_842));
FA_X1 i_415 (.CO (n_855), .S (n_854), .A (n_795), .B (n_793), .CI (n_791));
FA_X1 i_414 (.CO (n_853), .S (n_852), .A (n_787), .B (n_785), .CI (n_840));
FA_X1 i_413 (.CO (n_851), .S (n_850), .A (n_894), .B (n_937), .CI (n_789));
FA_X1 i_412 (.CO (n_849), .S (n_848), .A (n_783), .B (n_838), .CI (n_836));
FA_X1 i_411 (.CO (n_847), .S (n_846), .A (n_816), .B (n_814), .CI (n_812));
FA_X1 i_410 (.CO (n_845), .S (n_844), .A (n_822), .B (n_820), .CI (n_818));
FA_X1 i_409 (.CO (n_843), .S (n_842), .A (n_828), .B (n_826), .CI (n_824));
FA_X1 i_408 (.CO (n_841), .S (n_840), .A (n_779), .B (n_777), .CI (n_982));
FA_X1 i_407 (.CO (n_839), .S (n_838), .A (n_759), .B (n_757), .CI (n_781));
FA_X1 i_406 (.CO (n_829), .S (n_828), .A (n_2841), .B (n_2871), .CI (n_2899));
FA_X1 i_405 (.CO (n_827), .S (n_826), .A (n_2754), .B (n_2784), .CI (n_2812));
FA_X1 i_404 (.CO (n_825), .S (n_824), .A (n_2667), .B (n_2697), .CI (n_2725));
FA_X1 i_403 (.CO (n_823), .S (n_822), .A (n_2580), .B (n_2610), .CI (n_2638));
FA_X1 i_402 (.CO (n_821), .S (n_820), .A (n_2493), .B (n_2523), .CI (n_2551));
FA_X1 i_401 (.CO (n_819), .S (n_818), .A (n_2406), .B (n_2436), .CI (n_2464));
FA_X1 i_400 (.CO (n_817), .S (n_816), .A (n_2319), .B (n_2349), .CI (n_2377));
FA_X1 i_399 (.CO (n_815), .S (n_814), .A (n_2232), .B (n_2262), .CI (n_2290));
FA_X1 i_398 (.CO (n_813), .S (n_812), .A (n_2173), .B (n_2175), .CI (n_2203));
HA_X1 i_397 (.CO (n_811), .S (n_810), .A (n_753), .B (n_808));
FA_X1 i_396 (.CO (n_809), .S (n_808), .A (n_751), .B (n_804), .CI (n_806));
FA_X1 i_395 (.CO (n_807), .S (n_806), .A (n_800), .B (n_802), .CI (n_749));
FA_X1 i_394 (.CO (n_805), .S (n_804), .A (n_745), .B (n_747), .CI (n_798));
FA_X1 i_393 (.CO (n_803), .S (n_802), .A (n_792), .B (n_743), .CI (n_796));
FA_X1 i_392 (.CO (n_801), .S (n_800), .A (n_790), .B (n_741), .CI (n_794));
FA_X1 i_391 (.CO (n_799), .S (n_798), .A (n_788), .B (n_786), .CI (n_784));
FA_X1 i_390 (.CO (n_797), .S (n_796), .A (n_782), .B (n_739), .CI (n_737));
FA_X1 i_389 (.CO (n_795), .S (n_794), .A (n_733), .B (n_731), .CI (n_729));
FA_X1 i_388 (.CO (n_793), .S (n_792), .A (n_778), .B (n_776), .CI (n_735));
FA_X1 i_387 (.CO (n_791), .S (n_790), .A (n_756), .B (n_727), .CI (n_780));
FA_X1 i_386 (.CO (n_789), .S (n_788), .A (n_832), .B (n_834), .CI (n_758));
FA_X1 i_385 (.CO (n_787), .S (n_786), .A (n_884), .B (n_886), .CI (n_831));
FA_X1 i_384 (.CO (n_785), .S (n_784), .A (n_898), .B (n_900), .CI (n_870));
FA_X1 i_383 (.CO (n_783), .S (n_782), .A (n_725), .B (n_723), .CI (n_721));
FA_X1 i_382 (.CO (n_781), .S (n_780), .A (n_707), .B (n_705), .CI (n_703));
FA_X1 i_381 (.CO (n_779), .S (n_778), .A (n_713), .B (n_711), .CI (n_709));
FA_X1 i_380 (.CO (n_777), .S (n_776), .A (n_719), .B (n_717), .CI (n_715));
FA_X1 i_379 (.CO (n_759), .S (n_758), .A (n_2263), .B (n_2291), .CI (n_2320));
FA_X1 i_378 (.CO (n_757), .S (n_756), .A (n_2176), .B (n_2204), .CI (n_2233));
HA_X1 i_377 (.CO (n_755), .S (n_754), .A (n_699), .B (n_752));
FA_X1 i_376 (.CO (n_753), .S (n_752), .A (n_748), .B (n_697), .CI (n_750));
FA_X1 i_375 (.CO (n_751), .S (n_750), .A (n_744), .B (n_695), .CI (n_746));
FA_X1 i_374 (.CO (n_749), .S (n_748), .A (n_740), .B (n_693), .CI (n_742));
FA_X1 i_373 (.CO (n_747), .S (n_746), .A (n_736), .B (n_689), .CI (n_691));
FA_X1 i_372 (.CO (n_745), .S (n_744), .A (n_730), .B (n_687), .CI (n_738));
FA_X1 i_371 (.CO (n_743), .S (n_742), .A (n_683), .B (n_734), .CI (n_732));
FA_X1 i_370 (.CO (n_741), .S (n_740), .A (n_677), .B (n_728), .CI (n_685));
FA_X1 i_369 (.CO (n_739), .S (n_738), .A (n_722), .B (n_681), .CI (n_679));
FA_X1 i_368 (.CO (n_737), .S (n_736), .A (n_675), .B (n_726), .CI (n_724));
FA_X1 i_367 (.CO (n_735), .S (n_734), .A (n_706), .B (n_704), .CI (n_702));
FA_X1 i_366 (.CO (n_733), .S (n_732), .A (n_712), .B (n_710), .CI (n_708));
FA_X1 i_365 (.CO (n_731), .S (n_730), .A (n_718), .B (n_716), .CI (n_714));
FA_X1 i_364 (.CO (n_729), .S (n_728), .A (n_671), .B (n_669), .CI (n_720));
FA_X1 i_363 (.CO (n_727), .S (n_726), .A (n_653), .B (n_651), .CI (n_673));
FA_X1 i_362 (.CO (n_725), .S (n_724), .A (n_659), .B (n_657), .CI (n_655));
FA_X1 i_361 (.CO (n_723), .S (n_722), .A (n_665), .B (n_663), .CI (n_661));
FA_X1 i_360 (.CO (n_721), .S (n_720), .A (n_2988), .B (n_3016), .CI (n_667));
FA_X1 i_359 (.CO (n_719), .S (n_718), .A (n_2901), .B (n_2930), .CI (n_2959));
FA_X1 i_358 (.CO (n_717), .S (n_716), .A (n_2814), .B (n_2843), .CI (n_2873));
FA_X1 i_357 (.CO (n_715), .S (n_714), .A (n_2727), .B (n_2756), .CI (n_2786));
FA_X1 i_356 (.CO (n_713), .S (n_712), .A (n_2640), .B (n_2669), .CI (n_2699));
FA_X1 i_355 (.CO (n_711), .S (n_710), .A (n_2553), .B (n_2582), .CI (n_2612));
FA_X1 i_354 (.CO (n_709), .S (n_708), .A (n_2466), .B (n_2495), .CI (n_2525));
FA_X1 i_353 (.CO (n_707), .S (n_706), .A (n_2379), .B (n_2408), .CI (n_2438));
FA_X1 i_352 (.CO (n_705), .S (n_704), .A (n_2292), .B (n_2321), .CI (n_2351));
FA_X1 i_351 (.CO (n_703), .S (n_702), .A (n_2205), .B (n_2234), .CI (n_2264));
HA_X1 i_350 (.CO (n_701), .S (n_700), .A (n_647), .B (n_698));
FA_X1 i_349 (.CO (n_699), .S (n_698), .A (n_694), .B (n_645), .CI (n_696));
FA_X1 i_348 (.CO (n_697), .S (n_696), .A (n_690), .B (n_643), .CI (n_692));
FA_X1 i_347 (.CO (n_695), .S (n_694), .A (n_686), .B (n_688), .CI (n_641));
FA_X1 i_346 (.CO (n_693), .S (n_692), .A (n_684), .B (n_682), .CI (n_639));
FA_X1 i_345 (.CO (n_691), .S (n_690), .A (n_678), .B (n_676), .CI (n_637));
FA_X1 i_344 (.CO (n_689), .S (n_688), .A (n_635), .B (n_633), .CI (n_680));
FA_X1 i_343 (.CO (n_687), .S (n_686), .A (n_625), .B (n_631), .CI (n_674));
FA_X1 i_342 (.CO (n_685), .S (n_684), .A (n_668), .B (n_629), .CI (n_627));
FA_X1 i_341 (.CO (n_683), .S (n_682), .A (n_623), .B (n_672), .CI (n_670));
FA_X1 i_340 (.CO (n_681), .S (n_680), .A (n_654), .B (n_652), .CI (n_650));
FA_X1 i_339 (.CO (n_679), .S (n_678), .A (n_660), .B (n_658), .CI (n_656));
FA_X1 i_338 (.CO (n_677), .S (n_676), .A (n_666), .B (n_664), .CI (n_662));
FA_X1 i_337 (.CO (n_675), .S (n_674), .A (n_601), .B (n_621), .CI (n_619));
FA_X1 i_336 (.CO (n_673), .S (n_672), .A (n_607), .B (n_605), .CI (n_603));
FA_X1 i_335 (.CO (n_671), .S (n_670), .A (n_613), .B (n_611), .CI (n_609));
FA_X1 i_334 (.CO (n_669), .S (n_668), .A (n_3017), .B (n_617), .CI (n_615));
FA_X1 i_333 (.CO (n_667), .S (n_666), .A (n_2931), .B (n_2960), .CI (n_2989));
FA_X1 i_332 (.CO (n_665), .S (n_664), .A (n_2844), .B (n_2874), .CI (n_2902));
FA_X1 i_331 (.CO (n_663), .S (n_662), .A (n_2757), .B (n_2787), .CI (n_2815));
FA_X1 i_330 (.CO (n_661), .S (n_660), .A (n_2670), .B (n_2700), .CI (n_2728));
FA_X1 i_329 (.CO (n_659), .S (n_658), .A (n_2583), .B (n_2613), .CI (n_2641));
FA_X1 i_328 (.CO (n_657), .S (n_656), .A (n_2496), .B (n_2526), .CI (n_2554));
FA_X1 i_327 (.CO (n_655), .S (n_654), .A (n_2409), .B (n_2439), .CI (n_2467));
FA_X1 i_326 (.CO (n_653), .S (n_652), .A (n_2322), .B (n_2352), .CI (n_2380));
FA_X1 i_325 (.CO (n_651), .S (n_650), .A (n_2235), .B (n_2265), .CI (n_2293));
HA_X1 i_324 (.CO (n_649), .S (n_648), .A (n_597), .B (n_646));
FA_X1 i_323 (.CO (n_647), .S (n_646), .A (n_642), .B (n_595), .CI (n_644));
FA_X1 i_322 (.CO (n_645), .S (n_644), .A (n_638), .B (n_593), .CI (n_640));
FA_X1 i_321 (.CO (n_643), .S (n_642), .A (n_589), .B (n_636), .CI (n_591));
FA_X1 i_320 (.CO (n_641), .S (n_640), .A (n_587), .B (n_634), .CI (n_632));
FA_X1 i_319 (.CO (n_639), .S (n_638), .A (n_630), .B (n_628), .CI (n_626));
FA_X1 i_318 (.CO (n_637), .S (n_636), .A (n_624), .B (n_585), .CI (n_583));
FA_X1 i_317 (.CO (n_635), .S (n_634), .A (n_581), .B (n_579), .CI (n_577));
FA_X1 i_316 (.CO (n_633), .S (n_632), .A (n_622), .B (n_620), .CI (n_618));
FA_X1 i_315 (.CO (n_631), .S (n_630), .A (n_602), .B (n_600), .CI (n_575));
FA_X1 i_314 (.CO (n_629), .S (n_628), .A (n_608), .B (n_606), .CI (n_604));
FA_X1 i_313 (.CO (n_627), .S (n_626), .A (n_614), .B (n_612), .CI (n_610));
FA_X1 i_312 (.CO (n_625), .S (n_624), .A (n_571), .B (n_569), .CI (n_616));
FA_X1 i_311 (.CO (n_623), .S (n_622), .A (n_555), .B (n_553), .CI (n_573));
FA_X1 i_310 (.CO (n_621), .S (n_620), .A (n_561), .B (n_559), .CI (n_557));
FA_X1 i_309 (.CO (n_619), .S (n_618), .A (n_567), .B (n_565), .CI (n_563));
FA_X1 i_308 (.CO (n_617), .S (n_616), .A (n_2961), .B (n_2990), .CI (n_3018));
FA_X1 i_307 (.CO (n_615), .S (n_614), .A (n_2875), .B (n_2903), .CI (n_2932));
FA_X1 i_306 (.CO (n_613), .S (n_612), .A (n_2788), .B (n_2816), .CI (n_2845));
FA_X1 i_305 (.CO (n_611), .S (n_610), .A (n_2701), .B (n_2729), .CI (n_2758));
FA_X1 i_304 (.CO (n_609), .S (n_608), .A (n_2614), .B (n_2642), .CI (n_2671));
FA_X1 i_303 (.CO (n_607), .S (n_606), .A (n_2527), .B (n_2555), .CI (n_2584));
FA_X1 i_302 (.CO (n_605), .S (n_604), .A (n_2440), .B (n_2468), .CI (n_2497));
FA_X1 i_301 (.CO (n_603), .S (n_602), .A (n_2353), .B (n_2381), .CI (n_2410));
FA_X1 i_300 (.CO (n_601), .S (n_600), .A (n_2266), .B (n_2294), .CI (n_2323));
HA_X1 i_299 (.CO (n_599), .S (n_598), .A (n_549), .B (n_551));
FA_X1 i_298 (.CO (n_597), .S (n_596), .A (n_547), .B (n_592), .CI (n_594));
FA_X1 i_297 (.CO (n_595), .S (n_594), .A (n_545), .B (n_588), .CI (n_590));
FA_X1 i_296 (.CO (n_593), .S (n_592), .A (n_541), .B (n_586), .CI (n_543));
FA_X1 i_295 (.CO (n_591), .S (n_590), .A (n_539), .B (n_584), .CI (n_582));
FA_X1 i_294 (.CO (n_589), .S (n_588), .A (n_580), .B (n_578), .CI (n_576));
FA_X1 i_293 (.CO (n_587), .S (n_586), .A (n_574), .B (n_537), .CI (n_535));
FA_X1 i_292 (.CO (n_585), .S (n_584), .A (n_533), .B (n_531), .CI (n_529));
FA_X1 i_291 (.CO (n_583), .S (n_582), .A (n_552), .B (n_572), .CI (n_570));
FA_X1 i_290 (.CO (n_581), .S (n_580), .A (n_558), .B (n_556), .CI (n_554));
FA_X1 i_289 (.CO (n_579), .S (n_578), .A (n_564), .B (n_562), .CI (n_560));
FA_X1 i_288 (.CO (n_577), .S (n_576), .A (n_523), .B (n_568), .CI (n_566));
FA_X1 i_287 (.CO (n_575), .S (n_574), .A (n_507), .B (n_527), .CI (n_525));
FA_X1 i_286 (.CO (n_573), .S (n_572), .A (n_513), .B (n_511), .CI (n_509));
FA_X1 i_285 (.CO (n_571), .S (n_570), .A (n_519), .B (n_517), .CI (n_515));
FA_X1 i_284 (.CO (n_569), .S (n_568), .A (n_2991), .B (n_3019), .CI (n_521));
FA_X1 i_283 (.CO (n_567), .S (n_566), .A (n_2904), .B (n_2933), .CI (n_2962));
FA_X1 i_282 (.CO (n_565), .S (n_564), .A (n_2817), .B (n_2846), .CI (n_2876));
FA_X1 i_281 (.CO (n_563), .S (n_562), .A (n_2730), .B (n_2759), .CI (n_2789));
FA_X1 i_280 (.CO (n_561), .S (n_560), .A (n_2643), .B (n_2672), .CI (n_2702));
FA_X1 i_279 (.CO (n_559), .S (n_558), .A (n_2556), .B (n_2585), .CI (n_2615));
FA_X1 i_278 (.CO (n_557), .S (n_556), .A (n_2469), .B (n_2498), .CI (n_2528));
FA_X1 i_277 (.CO (n_555), .S (n_554), .A (n_2382), .B (n_2411), .CI (n_2441));
FA_X1 i_276 (.CO (n_553), .S (n_552), .A (n_2295), .B (n_2324), .CI (n_2354));
HA_X1 i_275 (.CO (n_551), .S (n_550), .A (n_503), .B (n_548));
FA_X1 i_274 (.CO (n_549), .S (n_548), .A (n_544), .B (n_501), .CI (n_546));
FA_X1 i_273 (.CO (n_547), .S (n_546), .A (n_499), .B (n_540), .CI (n_542));
FA_X1 i_272 (.CO (n_545), .S (n_544), .A (n_536), .B (n_495), .CI (n_497));
FA_X1 i_271 (.CO (n_543), .S (n_542), .A (n_534), .B (n_493), .CI (n_538));
FA_X1 i_270 (.CO (n_541), .S (n_540), .A (n_491), .B (n_532), .CI (n_530));
FA_X1 i_269 (.CO (n_539), .S (n_538), .A (n_487), .B (n_485), .CI (n_528));
FA_X1 i_268 (.CO (n_537), .S (n_536), .A (n_524), .B (n_522), .CI (n_489));
FA_X1 i_267 (.CO (n_535), .S (n_534), .A (n_506), .B (n_483), .CI (n_526));
FA_X1 i_266 (.CO (n_533), .S (n_532), .A (n_512), .B (n_510), .CI (n_508));
FA_X1 i_265 (.CO (n_531), .S (n_530), .A (n_518), .B (n_516), .CI (n_514));
FA_X1 i_264 (.CO (n_529), .S (n_528), .A (n_481), .B (n_479), .CI (n_520));
FA_X1 i_263 (.CO (n_527), .S (n_526), .A (n_467), .B (n_465), .CI (n_463));
FA_X1 i_262 (.CO (n_525), .S (n_524), .A (n_473), .B (n_471), .CI (n_469));
FA_X1 i_261 (.CO (n_523), .S (n_522), .A (n_3020), .B (n_477), .CI (n_475));
FA_X1 i_260 (.CO (n_521), .S (n_520), .A (n_2934), .B (n_2963), .CI (n_2992));
FA_X1 i_259 (.CO (n_519), .S (n_518), .A (n_2847), .B (n_2877), .CI (n_2905));
FA_X1 i_258 (.CO (n_517), .S (n_516), .A (n_2760), .B (n_2790), .CI (n_2818));
FA_X1 i_257 (.CO (n_515), .S (n_514), .A (n_2673), .B (n_2703), .CI (n_2731));
FA_X1 i_256 (.CO (n_513), .S (n_512), .A (n_2586), .B (n_2616), .CI (n_2644));
FA_X1 i_255 (.CO (n_511), .S (n_510), .A (n_2499), .B (n_2529), .CI (n_2557));
FA_X1 i_254 (.CO (n_509), .S (n_508), .A (n_2412), .B (n_2442), .CI (n_2470));
FA_X1 i_253 (.CO (n_507), .S (n_506), .A (n_2325), .B (n_2355), .CI (n_2383));
HA_X1 i_252 (.CO (n_505), .S (n_504), .A (n_459), .B (n_502));
FA_X1 i_251 (.CO (n_503), .S (n_502), .A (n_498), .B (n_457), .CI (n_500));
FA_X1 i_250 (.CO (n_501), .S (n_500), .A (n_494), .B (n_455), .CI (n_496));
FA_X1 i_249 (.CO (n_499), .S (n_498), .A (n_492), .B (n_490), .CI (n_453));
FA_X1 i_248 (.CO (n_497), .S (n_496), .A (n_486), .B (n_484), .CI (n_451));
FA_X1 i_247 (.CO (n_495), .S (n_494), .A (n_449), .B (n_447), .CI (n_488));
FA_X1 i_246 (.CO (n_493), .S (n_492), .A (n_443), .B (n_441), .CI (n_482));
FA_X1 i_245 (.CO (n_491), .S (n_490), .A (n_480), .B (n_478), .CI (n_445));
FA_X1 i_244 (.CO (n_489), .S (n_488), .A (n_466), .B (n_464), .CI (n_462));
FA_X1 i_243 (.CO (n_487), .S (n_486), .A (n_472), .B (n_470), .CI (n_468));
FA_X1 i_242 (.CO (n_485), .S (n_484), .A (n_435), .B (n_476), .CI (n_474));
FA_X1 i_241 (.CO (n_483), .S (n_482), .A (n_421), .B (n_439), .CI (n_437));
FA_X1 i_240 (.CO (n_481), .S (n_480), .A (n_427), .B (n_425), .CI (n_423));
FA_X1 i_239 (.CO (n_479), .S (n_478), .A (n_433), .B (n_431), .CI (n_429));
FA_X1 i_238 (.CO (n_477), .S (n_476), .A (n_2964), .B (n_2993), .CI (n_3021));
FA_X1 i_237 (.CO (n_475), .S (n_474), .A (n_2878), .B (n_2906), .CI (n_2935));
FA_X1 i_236 (.CO (n_473), .S (n_472), .A (n_2791), .B (n_2819), .CI (n_2848));
FA_X1 i_235 (.CO (n_471), .S (n_470), .A (n_2704), .B (n_2732), .CI (n_2761));
FA_X1 i_234 (.CO (n_469), .S (n_468), .A (n_2617), .B (n_2645), .CI (n_2674));
FA_X1 i_233 (.CO (n_467), .S (n_466), .A (n_2530), .B (n_2558), .CI (n_2587));
FA_X1 i_232 (.CO (n_465), .S (n_464), .A (n_2443), .B (n_2471), .CI (n_2500));
FA_X1 i_231 (.CO (n_463), .S (n_462), .A (n_2356), .B (n_2384), .CI (n_2413));
HA_X1 i_230 (.CO (n_461), .S (n_460), .A (n_417), .B (n_458));
FA_X1 i_229 (.CO (n_459), .S (n_458), .A (n_454), .B (n_415), .CI (n_456));
FA_X1 i_228 (.CO (n_457), .S (n_456), .A (n_450), .B (n_413), .CI (n_452));
FA_X1 i_227 (.CO (n_455), .S (n_454), .A (n_409), .B (n_448), .CI (n_411));
FA_X1 i_226 (.CO (n_453), .S (n_452), .A (n_444), .B (n_442), .CI (n_446));
FA_X1 i_225 (.CO (n_451), .S (n_450), .A (n_440), .B (n_407), .CI (n_405));
FA_X1 i_224 (.CO (n_449), .S (n_448), .A (n_436), .B (n_403), .CI (n_401));
FA_X1 i_223 (.CO (n_447), .S (n_446), .A (n_420), .B (n_399), .CI (n_438));
FA_X1 i_222 (.CO (n_445), .S (n_444), .A (n_426), .B (n_424), .CI (n_422));
FA_X1 i_221 (.CO (n_443), .S (n_442), .A (n_432), .B (n_430), .CI (n_428));
FA_X1 i_220 (.CO (n_441), .S (n_440), .A (n_397), .B (n_395), .CI (n_434));
FA_X1 i_219 (.CO (n_439), .S (n_438), .A (n_385), .B (n_383), .CI (n_381));
FA_X1 i_218 (.CO (n_437), .S (n_436), .A (n_391), .B (n_389), .CI (n_387));
FA_X1 i_217 (.CO (n_435), .S (n_434), .A (n_2994), .B (n_3022), .CI (n_393));
FA_X1 i_216 (.CO (n_433), .S (n_432), .A (n_2907), .B (n_2936), .CI (n_2965));
FA_X1 i_215 (.CO (n_431), .S (n_430), .A (n_2820), .B (n_2849), .CI (n_2879));
FA_X1 i_214 (.CO (n_429), .S (n_428), .A (n_2733), .B (n_2762), .CI (n_2792));
FA_X1 i_213 (.CO (n_427), .S (n_426), .A (n_2646), .B (n_2675), .CI (n_2705));
FA_X1 i_212 (.CO (n_425), .S (n_424), .A (n_2559), .B (n_2588), .CI (n_2618));
FA_X1 i_211 (.CO (n_423), .S (n_422), .A (n_2472), .B (n_2501), .CI (n_2531));
FA_X1 i_210 (.CO (n_421), .S (n_420), .A (n_2385), .B (n_2414), .CI (n_2444));
HA_X1 i_209 (.CO (n_419), .S (n_418), .A (n_377), .B (n_416));
FA_X1 i_208 (.CO (n_417), .S (n_416), .A (n_375), .B (n_412), .CI (n_414));
FA_X1 i_207 (.CO (n_415), .S (n_414), .A (n_371), .B (n_373), .CI (n_410));
FA_X1 i_206 (.CO (n_413), .S (n_412), .A (n_369), .B (n_408), .CI (n_406));
FA_X1 i_205 (.CO (n_411), .S (n_410), .A (n_404), .B (n_402), .CI (n_400));
FA_X1 i_204 (.CO (n_409), .S (n_408), .A (n_363), .B (n_361), .CI (n_367));
FA_X1 i_203 (.CO (n_407), .S (n_406), .A (n_396), .B (n_394), .CI (n_365));
FA_X1 i_202 (.CO (n_405), .S (n_404), .A (n_382), .B (n_380), .CI (n_398));
FA_X1 i_201 (.CO (n_403), .S (n_402), .A (n_388), .B (n_386), .CI (n_384));
FA_X1 i_200 (.CO (n_401), .S (n_400), .A (n_357), .B (n_392), .CI (n_390));
FA_X1 i_199 (.CO (n_399), .S (n_398), .A (n_345), .B (n_343), .CI (n_359));
FA_X1 i_198 (.CO (n_397), .S (n_396), .A (n_351), .B (n_349), .CI (n_347));
FA_X1 i_197 (.CO (n_395), .S (n_394), .A (n_3023), .B (n_355), .CI (n_353));
FA_X1 i_196 (.CO (n_393), .S (n_392), .A (n_2937), .B (n_2966), .CI (n_2995));
FA_X1 i_195 (.CO (n_391), .S (n_390), .A (n_2850), .B (n_2880), .CI (n_2908));
FA_X1 i_194 (.CO (n_389), .S (n_388), .A (n_2763), .B (n_2793), .CI (n_2821));
FA_X1 i_193 (.CO (n_387), .S (n_386), .A (n_2676), .B (n_2706), .CI (n_2734));
FA_X1 i_192 (.CO (n_385), .S (n_384), .A (n_2589), .B (n_2619), .CI (n_2647));
FA_X1 i_191 (.CO (n_383), .S (n_382), .A (n_2502), .B (n_2532), .CI (n_2560));
FA_X1 i_190 (.CO (n_381), .S (n_380), .A (n_2415), .B (n_2445), .CI (n_2473));
HA_X1 i_189 (.CO (n_379), .S (n_378), .A (n_339), .B (n_341));
FA_X1 i_188 (.CO (n_377), .S (n_376), .A (n_337), .B (n_372), .CI (n_374));
FA_X1 i_187 (.CO (n_375), .S (n_374), .A (n_333), .B (n_335), .CI (n_370));
FA_X1 i_186 (.CO (n_373), .S (n_372), .A (n_362), .B (n_368), .CI (n_366));
FA_X1 i_185 (.CO (n_371), .S (n_370), .A (n_331), .B (n_329), .CI (n_364));
FA_X1 i_184 (.CO (n_369), .S (n_368), .A (n_327), .B (n_325), .CI (n_360));
FA_X1 i_183 (.CO (n_367), .S (n_366), .A (n_323), .B (n_358), .CI (n_356));
FA_X1 i_182 (.CO (n_365), .S (n_364), .A (n_346), .B (n_344), .CI (n_342));
FA_X1 i_181 (.CO (n_363), .S (n_362), .A (n_352), .B (n_350), .CI (n_348));
FA_X1 i_180 (.CO (n_361), .S (n_360), .A (n_321), .B (n_319), .CI (n_354));
FA_X1 i_179 (.CO (n_359), .S (n_358), .A (n_311), .B (n_309), .CI (n_307));
FA_X1 i_178 (.CO (n_357), .S (n_356), .A (n_317), .B (n_315), .CI (n_313));
FA_X1 i_177 (.CO (n_355), .S (n_354), .A (n_2967), .B (n_2996), .CI (n_3024));
FA_X1 i_176 (.CO (n_353), .S (n_352), .A (n_2881), .B (n_2909), .CI (n_2938));
FA_X1 i_175 (.CO (n_351), .S (n_350), .A (n_2794), .B (n_2822), .CI (n_2851));
FA_X1 i_174 (.CO (n_349), .S (n_348), .A (n_2707), .B (n_2735), .CI (n_2764));
FA_X1 i_173 (.CO (n_347), .S (n_346), .A (n_2620), .B (n_2648), .CI (n_2677));
FA_X1 i_172 (.CO (n_345), .S (n_344), .A (n_2533), .B (n_2561), .CI (n_2590));
FA_X1 i_171 (.CO (n_343), .S (n_342), .A (n_2446), .B (n_2474), .CI (n_2503));
HA_X1 i_170 (.CO (n_341), .S (n_340), .A (n_303), .B (n_338));
FA_X1 i_169 (.CO (n_339), .S (n_338), .A (n_334), .B (n_301), .CI (n_336));
FA_X1 i_168 (.CO (n_337), .S (n_336), .A (n_330), .B (n_299), .CI (n_332));
FA_X1 i_167 (.CO (n_335), .S (n_334), .A (n_326), .B (n_324), .CI (n_297));
FA_X1 i_166 (.CO (n_333), .S (n_332), .A (n_293), .B (n_295), .CI (n_328));
FA_X1 i_165 (.CO (n_331), .S (n_330), .A (n_320), .B (n_291), .CI (n_289));
FA_X1 i_164 (.CO (n_329), .S (n_328), .A (n_308), .B (n_306), .CI (n_322));
FA_X1 i_163 (.CO (n_327), .S (n_326), .A (n_314), .B (n_312), .CI (n_310));
FA_X1 i_162 (.CO (n_325), .S (n_324), .A (n_285), .B (n_318), .CI (n_316));
FA_X1 i_161 (.CO (n_323), .S (n_322), .A (n_275), .B (n_273), .CI (n_287));
FA_X1 i_160 (.CO (n_321), .S (n_320), .A (n_281), .B (n_279), .CI (n_277));
FA_X1 i_159 (.CO (n_319), .S (n_318), .A (n_2997), .B (n_3025), .CI (n_283));
FA_X1 i_158 (.CO (n_317), .S (n_316), .A (n_2910), .B (n_2939), .CI (n_2968));
FA_X1 i_157 (.CO (n_315), .S (n_314), .A (n_2823), .B (n_2852), .CI (n_2882));
FA_X1 i_156 (.CO (n_313), .S (n_312), .A (n_2736), .B (n_2765), .CI (n_2795));
FA_X1 i_155 (.CO (n_311), .S (n_310), .A (n_2649), .B (n_2678), .CI (n_2708));
FA_X1 i_154 (.CO (n_309), .S (n_308), .A (n_2562), .B (n_2591), .CI (n_2621));
FA_X1 i_153 (.CO (n_307), .S (n_306), .A (n_2475), .B (n_2504), .CI (n_2534));
HA_X1 i_152 (.CO (n_305), .S (n_304), .A (n_269), .B (n_302));
FA_X1 i_151 (.CO (n_303), .S (n_302), .A (n_267), .B (n_298), .CI (n_300));
FA_X1 i_150 (.CO (n_301), .S (n_300), .A (n_294), .B (n_265), .CI (n_296));
FA_X1 i_149 (.CO (n_299), .S (n_298), .A (n_261), .B (n_292), .CI (n_290));
FA_X1 i_148 (.CO (n_297), .S (n_296), .A (n_257), .B (n_288), .CI (n_263));
FA_X1 i_147 (.CO (n_295), .S (n_294), .A (n_286), .B (n_284), .CI (n_259));
FA_X1 i_146 (.CO (n_293), .S (n_292), .A (n_274), .B (n_272), .CI (n_255));
FA_X1 i_145 (.CO (n_291), .S (n_290), .A (n_280), .B (n_278), .CI (n_276));
FA_X1 i_144 (.CO (n_289), .S (n_288), .A (n_241), .B (n_253), .CI (n_282));
FA_X1 i_143 (.CO (n_287), .S (n_286), .A (n_247), .B (n_245), .CI (n_243));
FA_X1 i_142 (.CO (n_285), .S (n_284), .A (n_3026), .B (n_251), .CI (n_249));
FA_X1 i_141 (.CO (n_283), .S (n_282), .A (n_2940), .B (n_2969), .CI (n_2998));
FA_X1 i_140 (.CO (n_281), .S (n_280), .A (n_2853), .B (n_2883), .CI (n_2911));
FA_X1 i_139 (.CO (n_279), .S (n_278), .A (n_2766), .B (n_2796), .CI (n_2824));
FA_X1 i_138 (.CO (n_277), .S (n_276), .A (n_2679), .B (n_2709), .CI (n_2737));
FA_X1 i_137 (.CO (n_275), .S (n_274), .A (n_2592), .B (n_2622), .CI (n_2650));
FA_X1 i_136 (.CO (n_273), .S (n_272), .A (n_2505), .B (n_2535), .CI (n_2563));
HA_X1 i_135 (.CO (n_271), .S (n_270), .A (n_237), .B (n_239));
FA_X1 i_134 (.CO (n_269), .S (n_268), .A (n_235), .B (n_264), .CI (n_266));
FA_X1 i_133 (.CO (n_267), .S (n_266), .A (n_260), .B (n_262), .CI (n_233));
FA_X1 i_132 (.CO (n_265), .S (n_264), .A (n_231), .B (n_258), .CI (n_256));
FA_X1 i_131 (.CO (n_263), .S (n_262), .A (n_252), .B (n_229), .CI (n_227));
FA_X1 i_130 (.CO (n_261), .S (n_260), .A (n_240), .B (n_225), .CI (n_254));
FA_X1 i_129 (.CO (n_259), .S (n_258), .A (n_246), .B (n_244), .CI (n_242));
FA_X1 i_128 (.CO (n_257), .S (n_256), .A (n_221), .B (n_250), .CI (n_248));
FA_X1 i_127 (.CO (n_255), .S (n_254), .A (n_213), .B (n_211), .CI (n_223));
FA_X1 i_126 (.CO (n_253), .S (n_252), .A (n_219), .B (n_217), .CI (n_215));
FA_X1 i_125 (.CO (n_251), .S (n_250), .A (n_2970), .B (n_2999), .CI (n_3027));
FA_X1 i_124 (.CO (n_249), .S (n_248), .A (n_2884), .B (n_2912), .CI (n_2941));
FA_X1 i_123 (.CO (n_247), .S (n_246), .A (n_2797), .B (n_2825), .CI (n_2854));
FA_X1 i_122 (.CO (n_245), .S (n_244), .A (n_2710), .B (n_2738), .CI (n_2767));
FA_X1 i_121 (.CO (n_243), .S (n_242), .A (n_2623), .B (n_2651), .CI (n_2680));
FA_X1 i_120 (.CO (n_241), .S (n_240), .A (n_2536), .B (n_2564), .CI (n_2593));
HA_X1 i_119 (.CO (n_239), .S (n_238), .A (n_207), .B (n_209));
FA_X1 i_118 (.CO (n_237), .S (n_236), .A (n_232), .B (n_205), .CI (n_234));
FA_X1 i_117 (.CO (n_235), .S (n_234), .A (n_226), .B (n_230), .CI (n_203));
FA_X1 i_116 (.CO (n_233), .S (n_232), .A (n_224), .B (n_201), .CI (n_228));
FA_X1 i_115 (.CO (n_231), .S (n_230), .A (n_222), .B (n_199), .CI (n_197));
FA_X1 i_114 (.CO (n_229), .S (n_228), .A (n_214), .B (n_212), .CI (n_210));
FA_X1 i_113 (.CO (n_227), .S (n_226), .A (n_220), .B (n_218), .CI (n_216));
FA_X1 i_112 (.CO (n_225), .S (n_224), .A (n_183), .B (n_195), .CI (n_193));
FA_X1 i_111 (.CO (n_223), .S (n_222), .A (n_189), .B (n_187), .CI (n_185));
FA_X1 i_110 (.CO (n_221), .S (n_220), .A (n_3000), .B (n_3028), .CI (n_191));
FA_X1 i_109 (.CO (n_219), .S (n_218), .A (n_2913), .B (n_2942), .CI (n_2971));
FA_X1 i_108 (.CO (n_217), .S (n_216), .A (n_2826), .B (n_2855), .CI (n_2885));
FA_X1 i_107 (.CO (n_215), .S (n_214), .A (n_2739), .B (n_2768), .CI (n_2798));
FA_X1 i_106 (.CO (n_213), .S (n_212), .A (n_2652), .B (n_2681), .CI (n_2711));
FA_X1 i_105 (.CO (n_211), .S (n_210), .A (n_2565), .B (n_2594), .CI (n_2624));
HA_X1 i_104 (.CO (n_209), .S (n_208), .A (n_179), .B (n_181));
FA_X1 i_103 (.CO (n_207), .S (n_206), .A (n_177), .B (n_202), .CI (n_204));
FA_X1 i_102 (.CO (n_205), .S (n_204), .A (n_196), .B (n_175), .CI (n_200));
FA_X1 i_101 (.CO (n_203), .S (n_202), .A (n_171), .B (n_173), .CI (n_198));
FA_X1 i_100 (.CO (n_201), .S (n_200), .A (n_169), .B (n_194), .CI (n_192));
FA_X1 i_99 (.CO (n_199), .S (n_198), .A (n_186), .B (n_184), .CI (n_182));
FA_X1 i_98 (.CO (n_197), .S (n_196), .A (n_167), .B (n_190), .CI (n_188));
FA_X1 i_97 (.CO (n_195), .S (n_194), .A (n_161), .B (n_159), .CI (n_157));
FA_X1 i_96 (.CO (n_193), .S (n_192), .A (n_3029), .B (n_165), .CI (n_163));
FA_X1 i_95 (.CO (n_191), .S (n_190), .A (n_2943), .B (n_2972), .CI (n_3001));
FA_X1 i_94 (.CO (n_189), .S (n_188), .A (n_2856), .B (n_2886), .CI (n_2914));
FA_X1 i_93 (.CO (n_187), .S (n_186), .A (n_2769), .B (n_2799), .CI (n_2827));
FA_X1 i_92 (.CO (n_185), .S (n_184), .A (n_2682), .B (n_2712), .CI (n_2740));
FA_X1 i_91 (.CO (n_183), .S (n_182), .A (n_2595), .B (n_2625), .CI (n_2653));
HA_X1 i_90 (.CO (n_181), .S (n_180), .A (n_153), .B (n_155));
FA_X1 i_89 (.CO (n_179), .S (n_178), .A (n_174), .B (n_151), .CI (n_176));
FA_X1 i_88 (.CO (n_177), .S (n_176), .A (n_149), .B (n_172), .CI (n_170));
FA_X1 i_87 (.CO (n_175), .S (n_174), .A (n_147), .B (n_145), .CI (n_168));
FA_X1 i_86 (.CO (n_173), .S (n_172), .A (n_158), .B (n_156), .CI (n_166));
FA_X1 i_85 (.CO (n_171), .S (n_170), .A (n_164), .B (n_162), .CI (n_160));
FA_X1 i_84 (.CO (n_169), .S (n_168), .A (n_133), .B (n_143), .CI (n_141));
FA_X1 i_83 (.CO (n_167), .S (n_166), .A (n_139), .B (n_137), .CI (n_135));
FA_X1 i_82 (.CO (n_165), .S (n_164), .A (n_2973), .B (n_3002), .CI (n_3030));
FA_X1 i_81 (.CO (n_163), .S (n_162), .A (n_2887), .B (n_2915), .CI (n_2944));
FA_X1 i_80 (.CO (n_161), .S (n_160), .A (n_2800), .B (n_2828), .CI (n_2857));
FA_X1 i_79 (.CO (n_159), .S (n_158), .A (n_2713), .B (n_2741), .CI (n_2770));
FA_X1 i_78 (.CO (n_157), .S (n_156), .A (n_2626), .B (n_2654), .CI (n_2683));
HA_X1 i_77 (.CO (n_155), .S (n_154), .A (n_150), .B (n_131));
FA_X1 i_76 (.CO (n_153), .S (n_152), .A (n_148), .B (n_127), .CI (n_129));
FA_X1 i_75 (.CO (n_151), .S (n_150), .A (n_125), .B (n_146), .CI (n_144));
FA_X1 i_74 (.CO (n_149), .S (n_148), .A (n_121), .B (n_142), .CI (n_123));
FA_X1 i_73 (.CO (n_147), .S (n_146), .A (n_136), .B (n_134), .CI (n_132));
FA_X1 i_72 (.CO (n_145), .S (n_144), .A (n_119), .B (n_140), .CI (n_138));
FA_X1 i_71 (.CO (n_143), .S (n_142), .A (n_115), .B (n_113), .CI (n_111));
FA_X1 i_70 (.CO (n_141), .S (n_140), .A (n_3003), .B (n_3031), .CI (n_117));
FA_X1 i_69 (.CO (n_139), .S (n_138), .A (n_2916), .B (n_2945), .CI (n_2974));
FA_X1 i_68 (.CO (n_137), .S (n_136), .A (n_2829), .B (n_2858), .CI (n_2888));
FA_X1 i_67 (.CO (n_135), .S (n_134), .A (n_2742), .B (n_2771), .CI (n_2801));
FA_X1 i_66 (.CO (n_133), .S (n_132), .A (n_2655), .B (n_2684), .CI (n_2714));
HA_X1 i_65 (.CO (n_131), .S (n_130), .A (n_107), .B (n_109));
FA_X1 i_64 (.CO (n_129), .S (n_128), .A (n_105), .B (n_124), .CI (n_126));
FA_X1 i_63 (.CO (n_127), .S (n_126), .A (n_101), .B (n_103), .CI (n_122));
FA_X1 i_62 (.CO (n_125), .S (n_124), .A (n_110), .B (n_120), .CI (n_118));
FA_X1 i_61 (.CO (n_123), .S (n_122), .A (n_116), .B (n_114), .CI (n_112));
FA_X1 i_60 (.CO (n_121), .S (n_120), .A (n_93), .B (n_91), .CI (n_99));
FA_X1 i_59 (.CO (n_119), .S (n_118), .A (n_3032), .B (n_97), .CI (n_95));
FA_X1 i_58 (.CO (n_117), .S (n_116), .A (n_2946), .B (n_2975), .CI (n_3004));
FA_X1 i_57 (.CO (n_115), .S (n_114), .A (n_2859), .B (n_2889), .CI (n_2917));
FA_X1 i_56 (.CO (n_113), .S (n_112), .A (n_2772), .B (n_2802), .CI (n_2830));
FA_X1 i_55 (.CO (n_111), .S (n_110), .A (n_2685), .B (n_2715), .CI (n_2743));
HA_X1 i_54 (.CO (n_109), .S (n_108), .A (n_89), .B (n_87));
FA_X1 i_53 (.CO (n_107), .S (n_106), .A (n_102), .B (n_100), .CI (n_104));
FA_X1 i_52 (.CO (n_105), .S (n_104), .A (n_98), .B (n_83), .CI (n_85));
FA_X1 i_51 (.CO (n_103), .S (n_102), .A (n_92), .B (n_90), .CI (n_81));
FA_X1 i_50 (.CO (n_101), .S (n_100), .A (n_79), .B (n_96), .CI (n_94));
FA_X1 i_49 (.CO (n_99), .S (n_98), .A (n_77), .B (n_75), .CI (n_73));
FA_X1 i_48 (.CO (n_97), .S (n_96), .A (n_2976), .B (n_3005), .CI (n_3033));
FA_X1 i_47 (.CO (n_95), .S (n_94), .A (n_2890), .B (n_2918), .CI (n_2947));
FA_X1 i_46 (.CO (n_93), .S (n_92), .A (n_2803), .B (n_2831), .CI (n_2860));
FA_X1 i_45 (.CO (n_91), .S (n_90), .A (n_2716), .B (n_2744), .CI (n_2773));
HA_X1 i_44 (.CO (n_89), .S (n_88), .A (n_71), .B (n_69));
FA_X1 i_43 (.CO (n_87), .S (n_86), .A (n_67), .B (n_82), .CI (n_84));
FA_X1 i_42 (.CO (n_85), .S (n_84), .A (n_72), .B (n_80), .CI (n_65));
FA_X1 i_41 (.CO (n_83), .S (n_82), .A (n_78), .B (n_76), .CI (n_74));
FA_X1 i_40 (.CO (n_81), .S (n_80), .A (n_59), .B (n_57), .CI (n_63));
FA_X1 i_39 (.CO (n_79), .S (n_78), .A (n_3006), .B (n_3034), .CI (n_61));
FA_X1 i_38 (.CO (n_77), .S (n_76), .A (n_2919), .B (n_2948), .CI (n_2977));
FA_X1 i_37 (.CO (n_75), .S (n_74), .A (n_2832), .B (n_2861), .CI (n_2891));
FA_X1 i_36 (.CO (n_73), .S (n_72), .A (n_2745), .B (n_2774), .CI (n_2804));
HA_X1 i_35 (.CO (n_71), .S (n_70), .A (n_55), .B (n_53));
FA_X1 i_34 (.CO (n_69), .S (n_68), .A (n_51), .B (n_64), .CI (n_66));
FA_X1 i_33 (.CO (n_67), .S (n_66), .A (n_56), .B (n_49), .CI (n_62));
FA_X1 i_32 (.CO (n_65), .S (n_64), .A (n_43), .B (n_60), .CI (n_58));
FA_X1 i_31 (.CO (n_63), .S (n_62), .A (n_3035), .B (n_47), .CI (n_45));
FA_X1 i_30 (.CO (n_61), .S (n_60), .A (n_2949), .B (n_2978), .CI (n_3007));
FA_X1 i_29 (.CO (n_59), .S (n_58), .A (n_2862), .B (n_2892), .CI (n_2920));
FA_X1 i_28 (.CO (n_57), .S (n_56), .A (n_2775), .B (n_2805), .CI (n_2833));
HA_X1 i_27 (.CO (n_55), .S (n_54), .A (n_39), .B (n_50));
FA_X1 i_26 (.CO (n_53), .S (n_52), .A (n_48), .B (n_37), .CI (n_41));
FA_X1 i_25 (.CO (n_51), .S (n_50), .A (n_46), .B (n_44), .CI (n_42));
FA_X1 i_24 (.CO (n_49), .S (n_48), .A (n_33), .B (n_31), .CI (n_35));
FA_X1 i_23 (.CO (n_47), .S (n_46), .A (n_2979), .B (n_3008), .CI (n_3036));
FA_X1 i_22 (.CO (n_45), .S (n_44), .A (n_2893), .B (n_2921), .CI (n_2950));
FA_X1 i_21 (.CO (n_43), .S (n_42), .A (n_2806), .B (n_2834), .CI (n_2863));
HA_X1 i_20 (.CO (n_41), .S (n_40), .A (n_36), .B (n_27));
FA_X1 i_19 (.CO (n_39), .S (n_38), .A (n_32), .B (n_30), .CI (n_29));
FA_X1 i_18 (.CO (n_37), .S (n_36), .A (n_21), .B (n_25), .CI (n_34));
FA_X1 i_17 (.CO (n_35), .S (n_34), .A (n_3009), .B (n_3037), .CI (n_23));
FA_X1 i_16 (.CO (n_33), .S (n_32), .A (n_2922), .B (n_2951), .CI (n_2980));
FA_X1 i_15 (.CO (n_31), .S (n_30), .A (n_2835), .B (n_2864), .CI (n_2894));
HA_X1 i_14 (.CO (n_29), .S (n_28), .A (n_19), .B (n_17));
FA_X1 i_13 (.CO (n_27), .S (n_26), .A (n_22), .B (n_20), .CI (n_24));
FA_X1 i_12 (.CO (n_25), .S (n_24), .A (n_3038), .B (n_15), .CI (n_13));
FA_X1 i_11 (.CO (n_23), .S (n_22), .A (n_2952), .B (n_2981), .CI (n_3010));
FA_X1 i_10 (.CO (n_21), .S (n_20), .A (n_2865), .B (n_2895), .CI (n_2923));
HA_X1 i_9 (.CO (n_19), .S (n_18), .A (n_12), .B (n_11));
FA_X1 i_8 (.CO (n_17), .S (n_16), .A (n_7), .B (n_9), .CI (n_14));
FA_X1 i_7 (.CO (n_15), .S (n_14), .A (n_2982), .B (n_3011), .CI (n_3039));
FA_X1 i_6 (.CO (n_13), .S (n_12), .A (n_2896), .B (n_2924), .CI (n_2953));
HA_X1 i_5 (.CO (n_11), .S (n_10), .A (n_3), .B (n_8));
FA_X1 i_4 (.CO (n_9), .S (n_8), .A (n_3012), .B (n_3040), .CI (n_5));
FA_X1 i_3 (.CO (n_7), .S (n_6), .A (n_2925), .B (n_2954), .CI (n_2983));
HA_X1 i_2 (.CO (n_5), .S (n_4), .A (n_3041), .B (n_1));
FA_X1 i_1 (.CO (n_3), .S (n_2), .A (n_2955), .B (n_2984), .CI (n_3013));
HA_X1 i_0 (.CO (n_1), .S (n_0), .A (n_2985), .B (n_3397));

endmodule //datapath

module multiplyTimes (inputA, inputB, result);

output [63:0] result;
input [31:0] inputA;
input [31:0] inputB;


datapath i_0 (.result ({result[63], result[62], result[61], result[60], result[59], 
    result[58], result[57], result[56], result[55], result[54], result[53], result[52], 
    result[51], result[50], result[49], result[48], result[47], result[46], result[45], 
    result[44], result[43], result[42], result[41], result[40], result[39], result[38], 
    result[37], result[36], result[35], result[34], result[33], result[32], result[31], 
    result[30], result[29], result[28], result[27], result[26], result[25], result[24], 
    result[23], result[22], result[21], result[20], result[19], result[18], result[17], 
    result[16], result[15], result[14], result[13], result[12], result[11], result[10], 
    result[9], result[8], result[7], result[6], result[5], result[4], result[3], 
    result[2], result[1], result[0]}), .inputA ({inputA[31], inputA[30], inputA[29], 
    inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], inputA[22], 
    inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], inputA[15], 
    inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], inputA[8], 
    inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], inputA[1], 
    inputA[0]}), .inputB ({inputB[31], inputB[30], inputB[29], inputB[28], inputB[27], 
    inputB[26], inputB[25], inputB[24], inputB[23], inputB[22], inputB[21], inputB[20], 
    inputB[19], inputB[18], inputB[17], inputB[16], inputB[15], inputB[14], inputB[13], 
    inputB[12], inputB[11], inputB[10], inputB[9], inputB[8], inputB[7], inputB[6], 
    inputB[5], inputB[4], inputB[3], inputB[2], inputB[1], inputB[0]}));

endmodule //multiplyTimes

module registerNbits__0_6 (clk_CTS_0_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_0;
wire drc_ipo_n6;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CLOCK_slh__n32;
wire CLOCK_slh__n33;
wire CLOCK_slh__n36;
wire CLOCK_slh__n37;
wire CLOCK_slh__n40;
wire CLOCK_slh__n41;
wire CLOCK_slh__n44;
wire CLOCK_slh__n45;
wire CLOCK_slh__n48;
wire CLOCK_slh__n50;
wire CLOCK_slh__n52;
wire CLOCK_slh__n54;
wire CLOCK_slh__n56;
wire CLOCK_slh__n58;
wire CLOCK_slh__n60;
wire CLOCK_slh__n62;
wire CLOCK_slh__n64;
wire CLOCK_slh__n66;
wire CLOCK_slh__n68;
wire CLOCK_slh__n70;
wire CLOCK_slh__n72;
wire CLOCK_slh__n74;
wire CLOCK_slh__n76;
wire CLOCK_slh__n78;
wire CLOCK_slh__n80;
wire CLOCK_slh__n82;
wire CLOCK_slh__n84;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n44), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n58), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n36), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n40), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n48), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n32), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n82), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n80), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n84), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n78), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n74), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n68), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n66), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n64), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n56), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n62), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n54), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n72), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n52), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n50), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n70), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n76), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n60), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n6), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
BUF_X2 drc_ipo_c3 (.Z (out[31]), .A (drc_ipo_n6));
CLKBUF_X1 CLOCK_slh__c10 (.Z (CLOCK_slh__n33), .A (CLOCK_slh__n32));
CLKBUF_X1 CLOCK_slh__c11 (.Z (n_28), .A (CLOCK_slh__n33));
CLKBUF_X1 CLOCK_slh__c14 (.Z (CLOCK_slh__n37), .A (CLOCK_slh__n36));
CLKBUF_X1 CLOCK_slh__c15 (.Z (n_31), .A (CLOCK_slh__n37));
CLKBUF_X1 CLOCK_slh__c18 (.Z (CLOCK_slh__n41), .A (CLOCK_slh__n40));
CLKBUF_X1 CLOCK_slh__c19 (.Z (n_30), .A (CLOCK_slh__n41));
CLKBUF_X1 CLOCK_slh__c22 (.Z (CLOCK_slh__n45), .A (CLOCK_slh__n44));
CLKBUF_X1 CLOCK_slh__c23 (.Z (n_33), .A (CLOCK_slh__n45));
CLKBUF_X1 CLOCK_slh__c26 (.Z (n_29), .A (CLOCK_slh__n48));
CLKBUF_X1 CLOCK_slh__c28 (.Z (n_5), .A (CLOCK_slh__n50));
CLKBUF_X1 CLOCK_slh__c30 (.Z (n_6), .A (CLOCK_slh__n52));
CLKBUF_X1 CLOCK_slh__c32 (.Z (n_8), .A (CLOCK_slh__n54));
CLKBUF_X1 CLOCK_slh__c34 (.Z (n_11), .A (CLOCK_slh__n56));
CLKBUF_X1 CLOCK_slh__c36 (.Z (n_32), .A (CLOCK_slh__n58));
CLKBUF_X1 CLOCK_slh__c38 (.Z (n_2), .A (CLOCK_slh__n60));
CLKBUF_X1 CLOCK_slh__c40 (.Z (n_9), .A (CLOCK_slh__n62));
CLKBUF_X1 CLOCK_slh__c42 (.Z (n_12), .A (CLOCK_slh__n64));
CLKBUF_X1 CLOCK_slh__c44 (.Z (n_13), .A (CLOCK_slh__n66));
CLKBUF_X1 CLOCK_slh__c46 (.Z (n_14), .A (CLOCK_slh__n68));
CLKBUF_X1 CLOCK_slh__c48 (.Z (n_4), .A (CLOCK_slh__n70));
CLKBUF_X1 CLOCK_slh__c50 (.Z (n_7), .A (CLOCK_slh__n72));
CLKBUF_X1 CLOCK_slh__c52 (.Z (n_15), .A (CLOCK_slh__n74));
CLKBUF_X1 CLOCK_slh__c54 (.Z (n_3), .A (CLOCK_slh__n76));
CLKBUF_X1 CLOCK_slh__c56 (.Z (n_16), .A (CLOCK_slh__n78));
CLKBUF_X1 CLOCK_slh__c58 (.Z (n_18), .A (CLOCK_slh__n80));
CLKBUF_X1 CLOCK_slh__c60 (.Z (n_20), .A (CLOCK_slh__n82));
CLKBUF_X1 CLOCK_slh__c62 (.Z (n_17), .A (CLOCK_slh__n84));

endmodule //registerNbits__0_6

module registerNbits__0_3 (clk_CTS_0_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_0;
wire drc_ipo_n4;
wire drc_ipo_n2;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_29;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X2 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_29), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_29), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_29), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_29), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_29), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_29), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_29), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_29), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_29), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_29), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_29), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_29), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_29), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_29), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_29), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_29), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_29), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_29), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_29), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_29), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_29), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_29), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_29), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_29), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_29), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_29), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_29), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_29), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_29), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_29), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (drc_ipo_n2), .CK (CTS_n_tid1_29), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n4), .CK (CTS_n_tid1_29), .D (n_33));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n_tid1_29), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
BUF_X1 drc_ipo_c1 (.Z (out[30]), .A (drc_ipo_n2));
BUF_X1 drc_ipo_c2 (.Z (out[31]), .A (drc_ipo_n4));

endmodule //registerNbits__0_3

module integrationMult (clk, reset, en, inputA, inputB, result);

output [63:0] result;
input clk;
input en;
input [31:0] inputA;
input [31:0] inputB;
input reset;
wire CTS_n_tid0_3;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire \outB_reg[31] ;
wire \outB_reg[30] ;
wire \outB_reg[29] ;
wire \outB_reg[28] ;
wire \outB_reg[27] ;
wire \outB_reg[26] ;
wire \outB_reg[25] ;
wire \outB_reg[24] ;
wire \outB_reg[23] ;
wire \outB_reg[22] ;
wire \outB_reg[21] ;
wire \outB_reg[20] ;
wire \outB_reg[19] ;
wire \outB_reg[18] ;
wire \outB_reg[17] ;
wire \outB_reg[16] ;
wire \outB_reg[15] ;
wire \outB_reg[14] ;
wire \outB_reg[13] ;
wire \outB_reg[12] ;
wire \outB_reg[11] ;
wire \outB_reg[10] ;
wire \outB_reg[9] ;
wire \outB_reg[8] ;
wire \outB_reg[7] ;
wire \outB_reg[6] ;
wire \outB_reg[5] ;
wire \outB_reg[4] ;
wire \outB_reg[3] ;
wire \outB_reg[2] ;
wire \outB_reg[1] ;
wire \outB_reg[0] ;
wire \outA_reg[31] ;
wire \outA_reg[30] ;
wire \outA_reg[29] ;
wire \outA_reg[28] ;
wire \outA_reg[27] ;
wire \outA_reg[26] ;
wire \outA_reg[25] ;
wire \outA_reg[24] ;
wire \outA_reg[23] ;
wire \outA_reg[22] ;
wire \outA_reg[21] ;
wire \outA_reg[20] ;
wire \outA_reg[19] ;
wire \outA_reg[18] ;
wire \outA_reg[17] ;
wire \outA_reg[16] ;
wire \outA_reg[15] ;
wire \outA_reg[14] ;
wire \outA_reg[13] ;
wire \outA_reg[12] ;
wire \outA_reg[11] ;
wire \outA_reg[10] ;
wire \outA_reg[9] ;
wire \outA_reg[8] ;
wire \outA_reg[7] ;
wire \outA_reg[6] ;
wire \outA_reg[5] ;
wire \outA_reg[4] ;
wire \outA_reg[3] ;
wire \outA_reg[2] ;
wire \outA_reg[1] ;
wire \outA_reg[0] ;
wire CTS_n_tid0_4;
wire CLOCK_n_tid0_89;


registerNbits outA (.out ({result[31], result[30], result[29], result[28], result[27], 
    result[26], result[25], result[24], result[23], result[22], result[21], result[20], 
    result[19], result[18], result[17], result[16], result[15], result[14], result[13], 
    result[12], result[11], result[10], result[9], result[8], result[7], result[6], 
    result[5], result[4], result[3], result[2], result[1], result[0]}), .en (en), .inp ({
    \outB_reg[31] , \outB_reg[30] , \outB_reg[29] , \outB_reg[28] , \outB_reg[27] , 
    \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , \outB_reg[23] , \outB_reg[22] , 
    \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , \outB_reg[18] , \outB_reg[17] , 
    \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , \outB_reg[13] , \outB_reg[12] , 
    \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , \outB_reg[8] , \outB_reg[7] , 
    \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , 
    \outB_reg[0] }), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_4));
registerNbits__0_9 outB (.out ({result[63], result[62], result[61], result[60], result[59], 
    result[58], result[57], result[56], result[55], result[54], result[53], result[52], 
    result[51], result[50], result[49], result[48], result[47], result[46], result[45], 
    result[44], result[43], result[42], result[41], result[40], result[39], result[38], 
    result[37], result[36], result[35], result[34], result[33], result[32]}), .clk_CTS_0_PP_0 (CTS_n_tid0_3)
    , .clk_CTS_0_PP_1 (CTS_n_tid0_4), .en (en), .inp ({\outA_reg[31] , \outA_reg[30] , 
    \outA_reg[29] , \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , 
    \outA_reg[24] , \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , 
    \outA_reg[19] , \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , 
    \outA_reg[14] , \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , 
    \outA_reg[9] , \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , 
    \outA_reg[3] , \outA_reg[2] , \outA_reg[1] , \outA_reg[0] }), .reset (reset), .clk_CTS_0_PP_2 (CLOCK_n_tid0_89));
multiplyTimes multiplier (.result ({\outA_reg[31] , \outA_reg[30] , \outA_reg[29] , 
    \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , \outA_reg[24] , 
    \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , \outA_reg[19] , 
    \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , \outA_reg[14] , 
    \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , \outA_reg[9] , 
    \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , 
    \outA_reg[2] , \outA_reg[1] , \outA_reg[0] , \outB_reg[31] , \outB_reg[30] , 
    \outB_reg[29] , \outB_reg[28] , \outB_reg[27] , \outB_reg[26] , \outB_reg[25] , 
    \outB_reg[24] , \outB_reg[23] , \outB_reg[22] , \outB_reg[21] , \outB_reg[20] , 
    \outB_reg[19] , \outB_reg[18] , \outB_reg[17] , \outB_reg[16] , \outB_reg[15] , 
    \outB_reg[14] , \outB_reg[13] , \outB_reg[12] , \outB_reg[11] , \outB_reg[10] , 
    \outB_reg[9] , \outB_reg[8] , \outB_reg[7] , \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , 
    \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , \outB_reg[0] }), .inputA ({\A_reg[31] , 
    \A_reg[30] , \A_reg[29] , \A_reg[28] , \A_reg[27] , \A_reg[26] , \A_reg[25] , 
    \A_reg[24] , \A_reg[23] , \A_reg[22] , \A_reg[21] , \A_reg[20] , \A_reg[19] , 
    \A_reg[18] , \A_reg[17] , \A_reg[16] , \A_reg[15] , \A_reg[14] , \A_reg[13] , 
    \A_reg[12] , \A_reg[11] , \A_reg[10] , \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , 
    \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , \A_reg[1] , \A_reg[0] }), .inputB ({
    \B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , \B_reg[26] , 
    \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , \B_reg[20] , 
    \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , \B_reg[14] , 
    \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , \B_reg[8] , \B_reg[7] , 
    \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] }));
registerNbits__0_6 regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , 
    \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , 
    \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , 
    \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , 
    \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .en (en), .inp ({inputB[31], inputB[30], 
    inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], inputB[24], inputB[23], 
    inputB[22], inputB[21], inputB[20], inputB[19], inputB[18], inputB[17], inputB[16], 
    inputB[15], inputB[14], inputB[13], inputB[12], inputB[11], inputB[10], inputB[9], 
    inputB[8], inputB[7], inputB[6], inputB[5], inputB[4], inputB[3], inputB[2], 
    inputB[1], inputB[0]}), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_4));
registerNbits__0_3 regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .en (en), .inp ({inputA[31], inputA[30], 
    inputA[29], inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], 
    inputA[22], inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], 
    inputA[15], inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], 
    inputA[8], inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], 
    inputA[1], inputA[0]}), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_3));
BUF_X4 CTS_L1_tid0__c1_tid0__c31 (.Z (CLOCK_n_tid0_89), .A (clk));

endmodule //integrationMult


