module empty (a,b,sum);
input a,b;
output sum;
assign sum = a+b;

endmodule
