/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Nov  5 15:42:38 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 4142605925 */

module datapath__0_66(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_67(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_66 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_68(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_69(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_68 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_70(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_71(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_70 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_72(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_73(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_72 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_74(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_75(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_74 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_76(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_77(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_76 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_78(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_79(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_78 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_80(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_81(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_80 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_82(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_83(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_82 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_84(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_85(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_84 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_86(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_87(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_86 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_88(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_89(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_88 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_90(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_91(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_90 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_92(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_93(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_92 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_94(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_95(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_94 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_96(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_97(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_96 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_98(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_99(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_98 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_100(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_101(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_100 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_102(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_103(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_102 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_104(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_105(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_104 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_106(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_107(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_106 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_108(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_109(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_108 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_110(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_111(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_110 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_112(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_113(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_112 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_114(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_115(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_114 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_116(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_117(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_116 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_118(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_119(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_118 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_120(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_121(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_120 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_122(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_123(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_122 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_124(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_125(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_124 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_126(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_127(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_126 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_2(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(1'b0), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_3(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_2 i_0 (.in2(in2), .c_in(), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_4(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_5(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_4 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_6(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_7(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_6 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_8(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_9(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_8 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_10(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_11(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_10 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_12(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_13(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_12 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_14(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_15(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_14 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_16(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_17(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_16 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_18(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_19(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_18 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_20(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_21(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_20 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_22(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_23(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_22 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_24(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_25(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_24 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_26(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_27(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_26 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_28(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_29(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_28 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_30(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_31(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_30 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_32(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_33(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_32 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_34(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_35(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_34 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_36(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_37(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_36 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_38(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_39(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_38 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_40(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_41(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_40 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_42(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_43(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_42 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_44(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_45(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_44 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_46(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_47(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_46 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_48(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_49(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_48 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_50(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_51(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_50 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_52(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_53(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_52 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_54(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_55(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_54 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_56(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_57(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_56 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_58(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_59(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_58 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_60(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_61(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_60 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_62(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(in2), .CO(p_0[1]), .S(p_0[0]));
endmodule

module Fulladder__0_63(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_62 i_0 (.in2(in2), .c_in(c_in), .in1(in1), .p_0({c_out, sum}));
endmodule

module datapath__0_64(in2, c_in, in1, p_0);
   input in2;
   input c_in;
   input in1;
   output [1:0]p_0;

   FA_X1 i_0 (.A(c_in), .B(in1), .CI(1'b0), .CO(n_0), .S(p_0[0]));
endmodule

module Fulladder__0_65(in1, in2, c_in, c_out, sum);
   input in1;
   input in2;
   input c_in;
   output c_out;
   output sum;

   datapath__0_64 i_0 (.in2(), .c_in(c_in), .in1(in1), .p_0({uc_0, sum}));
endmodule

module RippelCarryAdder(in1, in2, c_in, c_out, of, sum);
   input [31:0]in1;
   input [31:0]in2;
   input c_in;
   output c_out;
   output of;
   output [31:0]sum;

   wire [32:0]carrys;

   Fulladder__0_3 genblk1_0_FA (.in1(in1[0]), .in2(in2[0]), .c_in(), .c_out(
      carrys[1]), .sum(sum[0]));
   Fulladder__0_5 genblk1_1_FA (.in1(in1[1]), .in2(in2[1]), .c_in(carrys[1]), 
      .c_out(carrys[2]), .sum(sum[1]));
   Fulladder__0_7 genblk1_2_FA (.in1(in1[2]), .in2(in2[2]), .c_in(carrys[2]), 
      .c_out(carrys[3]), .sum(sum[2]));
   Fulladder__0_9 genblk1_3_FA (.in1(in1[3]), .in2(in2[3]), .c_in(carrys[3]), 
      .c_out(carrys[4]), .sum(sum[3]));
   Fulladder__0_11 genblk1_4_FA (.in1(in1[4]), .in2(in2[4]), .c_in(carrys[4]), 
      .c_out(carrys[5]), .sum(sum[4]));
   Fulladder__0_13 genblk1_5_FA (.in1(in1[5]), .in2(in2[5]), .c_in(carrys[5]), 
      .c_out(carrys[6]), .sum(sum[5]));
   Fulladder__0_15 genblk1_6_FA (.in1(in1[6]), .in2(in2[6]), .c_in(carrys[6]), 
      .c_out(carrys[7]), .sum(sum[6]));
   Fulladder__0_17 genblk1_7_FA (.in1(in1[7]), .in2(in2[7]), .c_in(carrys[7]), 
      .c_out(carrys[8]), .sum(sum[7]));
   Fulladder__0_19 genblk1_8_FA (.in1(in1[8]), .in2(in2[8]), .c_in(carrys[8]), 
      .c_out(carrys[9]), .sum(sum[8]));
   Fulladder__0_21 genblk1_9_FA (.in1(in1[9]), .in2(in2[9]), .c_in(carrys[9]), 
      .c_out(carrys[10]), .sum(sum[9]));
   Fulladder__0_23 genblk1_10_FA (.in1(in1[10]), .in2(in2[10]), .c_in(carrys[10]), 
      .c_out(carrys[11]), .sum(sum[10]));
   Fulladder__0_25 genblk1_11_FA (.in1(in1[11]), .in2(in2[11]), .c_in(carrys[11]), 
      .c_out(carrys[12]), .sum(sum[11]));
   Fulladder__0_27 genblk1_12_FA (.in1(in1[12]), .in2(in2[12]), .c_in(carrys[12]), 
      .c_out(carrys[13]), .sum(sum[12]));
   Fulladder__0_29 genblk1_13_FA (.in1(in1[13]), .in2(in2[13]), .c_in(carrys[13]), 
      .c_out(carrys[14]), .sum(sum[13]));
   Fulladder__0_31 genblk1_14_FA (.in1(in1[14]), .in2(in2[14]), .c_in(carrys[14]), 
      .c_out(carrys[15]), .sum(sum[14]));
   Fulladder__0_33 genblk1_15_FA (.in1(in1[15]), .in2(in2[15]), .c_in(carrys[15]), 
      .c_out(carrys[16]), .sum(sum[15]));
   Fulladder__0_35 genblk1_16_FA (.in1(in1[16]), .in2(in2[16]), .c_in(carrys[16]), 
      .c_out(carrys[17]), .sum(sum[16]));
   Fulladder__0_37 genblk1_17_FA (.in1(in1[17]), .in2(in2[17]), .c_in(carrys[17]), 
      .c_out(carrys[18]), .sum(sum[17]));
   Fulladder__0_39 genblk1_18_FA (.in1(in1[18]), .in2(in2[18]), .c_in(carrys[18]), 
      .c_out(carrys[19]), .sum(sum[18]));
   Fulladder__0_41 genblk1_19_FA (.in1(in1[19]), .in2(in2[19]), .c_in(carrys[19]), 
      .c_out(carrys[20]), .sum(sum[19]));
   Fulladder__0_43 genblk1_20_FA (.in1(in1[20]), .in2(in2[20]), .c_in(carrys[20]), 
      .c_out(carrys[21]), .sum(sum[20]));
   Fulladder__0_45 genblk1_21_FA (.in1(in1[21]), .in2(in2[21]), .c_in(carrys[21]), 
      .c_out(carrys[22]), .sum(sum[21]));
   Fulladder__0_47 genblk1_22_FA (.in1(in1[22]), .in2(in2[22]), .c_in(carrys[22]), 
      .c_out(carrys[23]), .sum(sum[22]));
   Fulladder__0_49 genblk1_23_FA (.in1(in1[23]), .in2(in2[23]), .c_in(carrys[23]), 
      .c_out(carrys[24]), .sum(sum[23]));
   Fulladder__0_51 genblk1_24_FA (.in1(in1[24]), .in2(in2[24]), .c_in(carrys[24]), 
      .c_out(carrys[25]), .sum(sum[24]));
   Fulladder__0_53 genblk1_25_FA (.in1(in1[25]), .in2(in2[25]), .c_in(carrys[25]), 
      .c_out(carrys[26]), .sum(sum[25]));
   Fulladder__0_55 genblk1_26_FA (.in1(in1[26]), .in2(in2[26]), .c_in(carrys[26]), 
      .c_out(carrys[27]), .sum(sum[26]));
   Fulladder__0_57 genblk1_27_FA (.in1(in1[27]), .in2(in2[27]), .c_in(carrys[27]), 
      .c_out(carrys[28]), .sum(sum[27]));
   Fulladder__0_59 genblk1_28_FA (.in1(in1[28]), .in2(in2[28]), .c_in(carrys[28]), 
      .c_out(carrys[29]), .sum(sum[28]));
   Fulladder__0_61 genblk1_29_FA (.in1(in1[29]), .in2(in2[29]), .c_in(carrys[29]), 
      .c_out(carrys[30]), .sum(sum[29]));
   Fulladder__0_63 genblk1_30_FA (.in1(in1[30]), .in2(in2[30]), .c_in(carrys[30]), 
      .c_out(carrys[31]), .sum(sum[30]));
   Fulladder__0_65 genblk1_31_FA (.in1(in1[31]), .in2(), .c_in(carrys[31]), 
      .c_out(), .sum(sum[31]));
endmodule

module overflow(A, B, sign, of);
   input A;
   input B;
   input sign;
   output of;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   INV_X1 i_0_0 (.A(B), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(A), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(sign), .ZN(n_0_2));
   OAI33_X1 i_0_3 (.A1(n_0_0), .A2(n_0_1), .A3(sign), .B1(n_0_2), .B2(A), 
      .B3(B), .ZN(of));
endmodule

module CarrySaveAdder(x, y, z, s, cout, of);
   input [31:0]x;
   input [31:0]y;
   input [31:0]z;
   output [31:0]s;
   output cout;
   output of;

   wire [31:0]r;
   wire [31:0]c;

   Fulladder__0_67 f31 (.in1(x[31]), .in2(y[31]), .c_in(z[31]), .c_out(c[31]), 
      .sum(r[31]));
   Fulladder__0_69 f30 (.in1(x[30]), .in2(y[30]), .c_in(z[30]), .c_out(c[30]), 
      .sum(r[30]));
   Fulladder__0_71 f29 (.in1(x[29]), .in2(y[29]), .c_in(z[29]), .c_out(c[29]), 
      .sum(r[29]));
   Fulladder__0_73 f28 (.in1(x[28]), .in2(y[28]), .c_in(z[28]), .c_out(c[28]), 
      .sum(r[28]));
   Fulladder__0_75 f27 (.in1(x[27]), .in2(y[27]), .c_in(z[27]), .c_out(c[27]), 
      .sum(r[27]));
   Fulladder__0_77 f26 (.in1(x[26]), .in2(y[26]), .c_in(z[26]), .c_out(c[26]), 
      .sum(r[26]));
   Fulladder__0_79 f25 (.in1(x[25]), .in2(y[25]), .c_in(z[25]), .c_out(c[25]), 
      .sum(r[25]));
   Fulladder__0_81 f24 (.in1(x[24]), .in2(y[24]), .c_in(z[24]), .c_out(c[24]), 
      .sum(r[24]));
   Fulladder__0_83 f23 (.in1(x[23]), .in2(y[23]), .c_in(z[23]), .c_out(c[23]), 
      .sum(r[23]));
   Fulladder__0_85 f22 (.in1(x[22]), .in2(y[22]), .c_in(z[22]), .c_out(c[22]), 
      .sum(r[22]));
   Fulladder__0_87 f21 (.in1(x[21]), .in2(y[21]), .c_in(z[21]), .c_out(c[21]), 
      .sum(r[21]));
   Fulladder__0_89 f20 (.in1(x[20]), .in2(y[20]), .c_in(z[20]), .c_out(c[20]), 
      .sum(r[20]));
   Fulladder__0_91 f19 (.in1(x[19]), .in2(y[19]), .c_in(z[19]), .c_out(c[19]), 
      .sum(r[19]));
   Fulladder__0_93 f18 (.in1(x[18]), .in2(y[18]), .c_in(z[18]), .c_out(c[18]), 
      .sum(r[18]));
   Fulladder__0_95 f17 (.in1(x[17]), .in2(y[17]), .c_in(z[17]), .c_out(c[17]), 
      .sum(r[17]));
   Fulladder__0_97 f16 (.in1(x[16]), .in2(y[16]), .c_in(z[16]), .c_out(c[16]), 
      .sum(r[16]));
   Fulladder__0_99 f15 (.in1(x[15]), .in2(y[15]), .c_in(z[15]), .c_out(c[15]), 
      .sum(r[15]));
   Fulladder__0_101 f14 (.in1(x[14]), .in2(y[14]), .c_in(z[14]), .c_out(c[14]), 
      .sum(r[14]));
   Fulladder__0_103 f13 (.in1(x[13]), .in2(y[13]), .c_in(z[13]), .c_out(c[13]), 
      .sum(r[13]));
   Fulladder__0_105 f12 (.in1(x[12]), .in2(y[12]), .c_in(z[12]), .c_out(c[12]), 
      .sum(r[12]));
   Fulladder__0_107 f11 (.in1(x[11]), .in2(y[11]), .c_in(z[11]), .c_out(c[11]), 
      .sum(r[11]));
   Fulladder__0_109 f10 (.in1(x[10]), .in2(y[10]), .c_in(z[10]), .c_out(c[10]), 
      .sum(r[10]));
   Fulladder__0_111 f9 (.in1(x[9]), .in2(y[9]), .c_in(z[9]), .c_out(c[9]), 
      .sum(r[9]));
   Fulladder__0_113 f8 (.in1(x[8]), .in2(y[8]), .c_in(z[8]), .c_out(c[8]), 
      .sum(r[8]));
   Fulladder__0_115 f7 (.in1(x[7]), .in2(y[7]), .c_in(z[7]), .c_out(c[7]), 
      .sum(r[7]));
   Fulladder__0_117 f6 (.in1(x[6]), .in2(y[6]), .c_in(z[6]), .c_out(c[6]), 
      .sum(r[6]));
   Fulladder__0_119 f5 (.in1(x[5]), .in2(y[5]), .c_in(z[5]), .c_out(c[5]), 
      .sum(r[5]));
   Fulladder__0_121 f4 (.in1(x[4]), .in2(y[4]), .c_in(z[4]), .c_out(c[4]), 
      .sum(r[4]));
   Fulladder__0_123 f3 (.in1(x[3]), .in2(y[3]), .c_in(z[3]), .c_out(c[3]), 
      .sum(r[3]));
   Fulladder__0_125 f2 (.in1(x[2]), .in2(y[2]), .c_in(z[2]), .c_out(c[2]), 
      .sum(r[2]));
   Fulladder__0_127 f1 (.in1(x[1]), .in2(y[1]), .c_in(z[1]), .c_out(c[1]), 
      .sum(r[1]));
   Fulladder f0 (.in1(x[0]), .in2(y[0]), .c_in(z[0]), .c_out(c[0]), .sum(s[0]));
   RippelCarryAdder rca (.in1(c), .in2({uc_0, r[31], r[30], r[29], r[28], r[27], 
      r[26], r[25], r[24], r[23], r[22], r[21], r[20], r[19], r[18], r[17], 
      r[16], r[15], r[14], r[13], r[12], r[11], r[10], r[9], r[8], r[7], r[6], 
      r[5], r[4], r[3], r[2], r[1]}), .c_in(), .c_out(), .of(), .sum({cout, 
      s[31], s[30], s[29], s[28], s[27], s[26], s[25], s[24], s[23], s[22], 
      s[21], s[20], s[19], s[18], s[17], s[16], s[15], s[14], s[13], s[12], 
      s[11], s[10], s[9], s[8], s[7], s[6], s[5], s[4], s[3], s[2], s[1]}));
   overflow overFlow (.A(x[31]), .B(y[31]), .sign(s[31]), .of(of));
endmodule
