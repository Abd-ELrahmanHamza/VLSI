/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Jan  3 03:38:00 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3358275526 */

module registerNbits__0_84(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits__0_87(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module datapath(firstInputComplement, a);
   output [31:0]firstInputComplement;
   input [31:0]a;

   XOR2_X1 i_0 (.A(a[1]), .B(a[0]), .Z(firstInputComplement[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(firstInputComplement[2]));
   OAI21_X1 i_2 (.A(a[2]), .B1(a[1]), .B2(a[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(a[3]), .B(n_29), .Z(firstInputComplement[3]));
   XOR2_X1 i_4 (.A(a[4]), .B(n_28), .Z(firstInputComplement[4]));
   XOR2_X1 i_5 (.A(a[5]), .B(n_27), .Z(firstInputComplement[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(firstInputComplement[6]));
   OAI21_X1 i_7 (.A(a[6]), .B1(n_27), .B2(a[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(a[7]), .B(n_26), .Z(firstInputComplement[7]));
   XOR2_X1 i_9 (.A(a[8]), .B(n_25), .Z(firstInputComplement[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(firstInputComplement[9]));
   OAI21_X1 i_11 (.A(a[9]), .B1(n_25), .B2(a[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(a[10]), .B(n_24), .Z(firstInputComplement[10]));
   XNOR2_X1 i_13 (.A(a[11]), .B(n_23), .ZN(firstInputComplement[11]));
   XOR2_X1 i_14 (.A(a[12]), .B(n_22), .Z(firstInputComplement[12]));
   XNOR2_X1 i_15 (.A(a[13]), .B(n_21), .ZN(firstInputComplement[13]));
   XNOR2_X1 i_16 (.A(a[14]), .B(n_20), .ZN(firstInputComplement[14]));
   XOR2_X1 i_17 (.A(a[15]), .B(n_19), .Z(firstInputComplement[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(firstInputComplement[16]));
   OAI21_X1 i_19 (.A(a[16]), .B1(n_19), .B2(a[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(a[17]), .B(n_18), .Z(firstInputComplement[17]));
   XOR2_X1 i_21 (.A(a[18]), .B(n_17), .Z(firstInputComplement[18]));
   XNOR2_X1 i_22 (.A(a[19]), .B(n_16), .ZN(firstInputComplement[19]));
   XNOR2_X1 i_23 (.A(a[20]), .B(n_15), .ZN(firstInputComplement[20]));
   XNOR2_X1 i_24 (.A(a[21]), .B(n_14), .ZN(firstInputComplement[21]));
   XOR2_X1 i_25 (.A(a[22]), .B(n_13), .Z(firstInputComplement[22]));
   XOR2_X1 i_26 (.A(a[23]), .B(n_12), .Z(firstInputComplement[23]));
   XNOR2_X1 i_27 (.A(a[24]), .B(n_11), .ZN(firstInputComplement[24]));
   XNOR2_X1 i_28 (.A(a[25]), .B(n_10), .ZN(firstInputComplement[25]));
   XOR2_X1 i_29 (.A(a[26]), .B(n_9), .Z(firstInputComplement[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(firstInputComplement[27]));
   OAI21_X1 i_31 (.A(a[27]), .B1(n_9), .B2(a[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(a[28]), .B(n_8), .Z(firstInputComplement[28]));
   XNOR2_X1 i_33 (.A(a[29]), .B(n_7), .ZN(firstInputComplement[29]));
   XNOR2_X1 i_34 (.A(a[30]), .B(n_6), .ZN(firstInputComplement[30]));
   XNOR2_X1 i_35 (.A(a[31]), .B(n_5), .ZN(firstInputComplement[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(a[28]), .A3(a[29]), .A4(a[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(a[28]), .A3(a[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(a[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(a[26]), .A3(a[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(a[23]), .A3(a[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(a[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(a[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(a[18]), .A3(a[19]), .A4(a[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(a[18]), .A3(a[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(a[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(a[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(a[15]), .A3(a[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(a[12]), .A3(a[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(a[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(a[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(a[8]), .A3(a[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(a[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(a[5]), .A3(a[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(a[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(a[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(a[2]), .A2(a[1]), .A3(a[0]), .ZN(n_29));
   INV_X1 i_61 (.A(a[11]), .ZN(n_30));
   INV_X1 i_62 (.A(a[14]), .ZN(n_31));
   INV_X1 i_63 (.A(a[21]), .ZN(n_32));
   INV_X1 i_64 (.A(a[25]), .ZN(n_33));
endmodule

module datapath__0_74(p_0, aux, p_1);
   input [63:0]p_0;
   input [63:0]aux;
   output [63:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_366), .B1(p_0[0]), .B2(aux[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_366), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_365), .B1(p_0[1]), .B2(aux[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_364), .B(n_2), .ZN(p_1[2]));
   OAI21_X1 i_5 (.A(n_369), .B1(p_0[2]), .B2(aux[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_363), .B(n_3), .Z(p_1[3]));
   OAI21_X1 i_7 (.A(n_370), .B1(n_376), .B2(n_372), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_361), .B(n_10), .Z(p_1[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_358), .A2(n_349), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(aux[6]), .B1(n_349), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_359), .B1(p_0[5]), .B2(aux[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_359), .B1(n_353), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_356), .B1(n_361), .B2(n_354), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_354), .B1(p_0[4]), .B2(aux[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_360), .A2(n_351), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_347), .B(n_18), .ZN(p_1[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_1[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_344), .A2(n_335), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(aux[10]), .B1(n_335), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_345), .B1(p_0[9]), .B2(aux[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_345), .B1(n_339), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_342), .B1(n_347), .B2(n_340), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_342), .B1(p_0[8]), .B2(aux[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_346), .A2(n_337), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_333), .B(n_26), .Z(p_1[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_1[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_1[14]));
   NOR2_X1 i_35 (.A1(n_330), .A2(n_321), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_1[15]));
   OAI22_X1 i_37 (.A1(p_0[14]), .A2(aux[14]), .B1(n_321), .B2(n_23), .ZN(n_21));
   AOI21_X1 i_38 (.A(n_331), .B1(p_0[13]), .B2(aux[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_331), .B1(n_325), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_328), .B1(n_333), .B2(n_326), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_326), .B1(p_0[12]), .B2(aux[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_332), .A2(n_323), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_319), .B(n_34), .Z(p_1[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_1[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_1[18]));
   NOR2_X1 i_47 (.A1(n_285), .A2(n_275), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_1[19]));
   OAI21_X1 i_49 (.A(n_284), .B1(n_275), .B2(n_31), .ZN(n_29));
   NOR2_X1 i_50 (.A1(n_287), .A2(n_277), .ZN(n_30));
   INV_X1 i_51 (.A(n_32), .ZN(n_31));
   OAI21_X1 i_52 (.A(n_286), .B1(n_277), .B2(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_282), .B1(n_319), .B2(n_279), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_279), .B1(p_0[16]), .B2(aux[16]), .ZN(n_34));
   AOI21_X1 i_55 (.A(n_289), .B1(p_0[19]), .B2(aux[19]), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_63), .B(n_42), .Z(p_1[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_1[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_1[22]));
   NOR2_X1 i_59 (.A1(n_313), .A2(n_257), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_1[23]));
   OAI21_X1 i_61 (.A(n_312), .B1(n_257), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_315), .A2(n_259), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_314), .B1(n_259), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_318), .B1(n_261), .B2(n_63), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_261), .B1(p_0[20]), .B2(aux[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_317), .B1(p_0[23]), .B2(aux[23]), .ZN(n_43));
   XOR2_X1 i_68 (.A(n_61), .B(n_50), .Z(p_1[24]));
   XOR2_X1 i_69 (.A(n_49), .B(n_46), .Z(p_1[25]));
   XOR2_X1 i_70 (.A(n_47), .B(n_44), .Z(p_1[26]));
   NOR2_X1 i_71 (.A1(n_296), .A2(n_269), .ZN(n_44));
   XNOR2_X1 i_72 (.A(n_51), .B(n_45), .ZN(p_1[27]));
   OAI21_X1 i_73 (.A(n_295), .B1(n_269), .B2(n_47), .ZN(n_45));
   NOR2_X1 i_74 (.A1(n_298), .A2(n_271), .ZN(n_46));
   INV_X1 i_75 (.A(n_48), .ZN(n_47));
   OAI21_X1 i_76 (.A(n_297), .B1(n_271), .B2(n_49), .ZN(n_48));
   AOI21_X1 i_77 (.A(n_293), .B1(n_273), .B2(n_61), .ZN(n_49));
   OAI21_X1 i_78 (.A(n_273), .B1(p_0[24]), .B2(aux[24]), .ZN(n_50));
   AOI21_X1 i_79 (.A(n_300), .B1(p_0[27]), .B2(aux[27]), .ZN(n_51));
   XOR2_X1 i_80 (.A(n_59), .B(n_58), .Z(p_1[28]));
   XOR2_X1 i_81 (.A(n_57), .B(n_54), .Z(p_1[29]));
   XOR2_X1 i_82 (.A(n_55), .B(n_52), .Z(p_1[30]));
   NOR2_X1 i_83 (.A1(n_305), .A2(n_263), .ZN(n_52));
   XOR2_X1 i_84 (.A(n_65), .B(n_53), .Z(p_1[31]));
   OAI21_X1 i_85 (.A(n_304), .B1(n_263), .B2(n_55), .ZN(n_53));
   NOR2_X1 i_86 (.A1(n_307), .A2(n_266), .ZN(n_54));
   INV_X1 i_87 (.A(n_56), .ZN(n_55));
   OAI21_X1 i_88 (.A(n_306), .B1(n_266), .B2(n_57), .ZN(n_56));
   AOI21_X1 i_89 (.A(n_302), .B1(n_267), .B2(n_59), .ZN(n_57));
   OAI21_X1 i_90 (.A(n_267), .B1(p_0[28]), .B2(aux[28]), .ZN(n_58));
   INV_X1 i_91 (.A(n_60), .ZN(n_59));
   OAI21_X1 i_92 (.A(n_268), .B1(n_292), .B2(n_61), .ZN(n_60));
   INV_X1 i_93 (.A(n_62), .ZN(n_61));
   OAI21_X1 i_94 (.A(n_256), .B1(n_310), .B2(n_63), .ZN(n_62));
   INV_X1 i_95 (.A(n_64), .ZN(n_63));
   OAI21_X1 i_96 (.A(n_274), .B1(n_319), .B2(n_281), .ZN(n_64));
   OAI21_X1 i_97 (.A(n_308), .B1(n_377), .B2(n_373), .ZN(n_65));
   XOR2_X1 i_98 (.A(n_254), .B(n_72), .Z(p_1[32]));
   XOR2_X1 i_99 (.A(n_71), .B(n_68), .Z(p_1[33]));
   XOR2_X1 i_100 (.A(n_69), .B(n_66), .Z(p_1[34]));
   NOR2_X1 i_101 (.A1(n_223), .A2(n_213), .ZN(n_66));
   XNOR2_X1 i_102 (.A(n_73), .B(n_67), .ZN(p_1[35]));
   OAI21_X1 i_103 (.A(n_222), .B1(n_213), .B2(n_69), .ZN(n_67));
   NOR2_X1 i_104 (.A1(n_225), .A2(n_215), .ZN(n_68));
   INV_X1 i_105 (.A(n_70), .ZN(n_69));
   OAI21_X1 i_106 (.A(n_224), .B1(n_215), .B2(n_71), .ZN(n_70));
   AOI21_X1 i_107 (.A(n_220), .B1(n_254), .B2(n_217), .ZN(n_71));
   OAI21_X1 i_108 (.A(n_217), .B1(p_0[32]), .B2(aux[32]), .ZN(n_72));
   AOI21_X1 i_109 (.A(n_227), .B1(p_0[35]), .B2(aux[35]), .ZN(n_73));
   XOR2_X1 i_110 (.A(n_101), .B(n_80), .Z(p_1[36]));
   XOR2_X1 i_111 (.A(n_79), .B(n_76), .Z(p_1[37]));
   XOR2_X1 i_112 (.A(n_77), .B(n_74), .Z(p_1[38]));
   NOR2_X1 i_113 (.A1(n_248), .A2(n_206), .ZN(n_74));
   XNOR2_X1 i_114 (.A(n_81), .B(n_75), .ZN(p_1[39]));
   OAI21_X1 i_115 (.A(n_247), .B1(n_206), .B2(n_77), .ZN(n_75));
   NOR2_X1 i_116 (.A1(n_250), .A2(n_208), .ZN(n_76));
   INV_X1 i_117 (.A(n_78), .ZN(n_77));
   OAI21_X1 i_118 (.A(n_249), .B1(n_208), .B2(n_79), .ZN(n_78));
   AOI21_X1 i_119 (.A(n_253), .B1(n_210), .B2(n_101), .ZN(n_79));
   OAI21_X1 i_120 (.A(n_210), .B1(p_0[36]), .B2(aux[36]), .ZN(n_80));
   AOI21_X1 i_121 (.A(n_252), .B1(p_0[39]), .B2(aux[39]), .ZN(n_81));
   XOR2_X1 i_122 (.A(n_99), .B(n_88), .Z(p_1[40]));
   XOR2_X1 i_123 (.A(n_87), .B(n_84), .Z(p_1[41]));
   XOR2_X1 i_124 (.A(n_85), .B(n_82), .Z(p_1[42]));
   NOR2_X1 i_125 (.A1(n_234), .A2(n_192), .ZN(n_82));
   XNOR2_X1 i_126 (.A(n_89), .B(n_83), .ZN(p_1[43]));
   OAI21_X1 i_127 (.A(n_233), .B1(n_192), .B2(n_85), .ZN(n_83));
   NOR2_X1 i_128 (.A1(n_236), .A2(n_194), .ZN(n_84));
   INV_X1 i_129 (.A(n_86), .ZN(n_85));
   OAI21_X1 i_130 (.A(n_235), .B1(n_194), .B2(n_87), .ZN(n_86));
   AOI21_X1 i_131 (.A(n_231), .B1(n_196), .B2(n_99), .ZN(n_87));
   OAI21_X1 i_132 (.A(n_196), .B1(p_0[40]), .B2(aux[40]), .ZN(n_88));
   AOI21_X1 i_133 (.A(n_238), .B1(p_0[43]), .B2(aux[43]), .ZN(n_89));
   XNOR2_X1 i_134 (.A(n_98), .B(n_97), .ZN(p_1[44]));
   XOR2_X1 i_135 (.A(n_95), .B(n_94), .Z(p_1[45]));
   XNOR2_X1 i_136 (.A(n_91), .B(n_90), .ZN(p_1[46]));
   OAI22_X1 i_137 (.A1(p_0[45]), .A2(aux[45]), .B1(n_202), .B2(n_95), .ZN(n_90));
   NOR2_X1 i_138 (.A1(n_242), .A2(n_199), .ZN(n_91));
   XNOR2_X1 i_139 (.A(n_103), .B(n_92), .ZN(p_1[47]));
   OAI21_X1 i_140 (.A(n_93), .B1(n_241), .B2(n_199), .ZN(n_92));
   NAND3_X1 i_141 (.A1(n_200), .A2(n_94), .A3(n_96), .ZN(n_93));
   NOR2_X1 i_142 (.A1(n_243), .A2(n_202), .ZN(n_94));
   INV_X1 i_143 (.A(n_96), .ZN(n_95));
   OAI22_X1 i_144 (.A1(p_0[44]), .A2(aux[44]), .B1(n_203), .B2(n_98), .ZN(n_96));
   OAI21_X1 i_145 (.A(n_204), .B1(p_0[44]), .B2(aux[44]), .ZN(n_97));
   OAI21_X1 i_146 (.A(n_191), .B1(n_230), .B2(n_99), .ZN(n_98));
   INV_X1 i_147 (.A(n_100), .ZN(n_99));
   OAI21_X1 i_148 (.A(n_205), .B1(n_245), .B2(n_101), .ZN(n_100));
   INV_X1 i_149 (.A(n_102), .ZN(n_101));
   OAI21_X1 i_150 (.A(n_212), .B1(n_254), .B2(n_219), .ZN(n_102));
   AOI21_X1 i_151 (.A(n_244), .B1(p_0[47]), .B2(aux[47]), .ZN(n_103));
   XOR2_X1 i_152 (.A(n_189), .B(n_110), .Z(p_1[48]));
   XOR2_X1 i_153 (.A(n_109), .B(n_106), .Z(p_1[49]));
   XOR2_X1 i_154 (.A(n_107), .B(n_104), .Z(p_1[50]));
   NOR2_X1 i_155 (.A1(n_186), .A2(n_177), .ZN(n_104));
   XNOR2_X1 i_156 (.A(n_111), .B(n_105), .ZN(p_1[51]));
   OAI22_X1 i_157 (.A1(p_0[50]), .A2(aux[50]), .B1(n_177), .B2(n_107), .ZN(n_105));
   AOI21_X1 i_158 (.A(n_187), .B1(p_0[49]), .B2(aux[49]), .ZN(n_106));
   AOI21_X1 i_159 (.A(n_187), .B1(n_181), .B2(n_108), .ZN(n_107));
   INV_X1 i_160 (.A(n_109), .ZN(n_108));
   AOI21_X1 i_161 (.A(n_184), .B1(n_189), .B2(n_182), .ZN(n_109));
   OAI21_X1 i_162 (.A(n_182), .B1(p_0[48]), .B2(aux[48]), .ZN(n_110));
   NOR2_X1 i_163 (.A1(n_188), .A2(n_179), .ZN(n_111));
   XOR2_X1 i_164 (.A(n_175), .B(n_118), .Z(p_1[52]));
   XOR2_X1 i_165 (.A(n_117), .B(n_114), .Z(p_1[53]));
   XOR2_X1 i_166 (.A(n_115), .B(n_112), .Z(p_1[54]));
   NOR2_X1 i_167 (.A1(n_164), .A2(n_154), .ZN(n_112));
   XNOR2_X1 i_168 (.A(n_119), .B(n_113), .ZN(p_1[55]));
   OAI21_X1 i_169 (.A(n_163), .B1(n_154), .B2(n_115), .ZN(n_113));
   NOR2_X1 i_170 (.A1(n_166), .A2(n_156), .ZN(n_114));
   INV_X1 i_171 (.A(n_116), .ZN(n_115));
   OAI21_X1 i_172 (.A(n_165), .B1(n_156), .B2(n_117), .ZN(n_116));
   AOI21_X1 i_173 (.A(n_161), .B1(n_175), .B2(n_158), .ZN(n_117));
   OAI21_X1 i_174 (.A(n_158), .B1(p_0[52]), .B2(aux[52]), .ZN(n_118));
   AOI21_X1 i_175 (.A(n_168), .B1(p_0[55]), .B2(aux[55]), .ZN(n_119));
   XNOR2_X1 i_176 (.A(n_128), .B(n_127), .ZN(p_1[56]));
   XOR2_X1 i_177 (.A(n_125), .B(n_124), .Z(p_1[57]));
   XNOR2_X1 i_178 (.A(n_121), .B(n_120), .ZN(p_1[58]));
   OAI22_X1 i_179 (.A1(p_0[57]), .A2(aux[57]), .B1(n_149), .B2(n_125), .ZN(n_120));
   NOR2_X1 i_180 (.A1(n_172), .A2(n_145), .ZN(n_121));
   XNOR2_X1 i_181 (.A(n_129), .B(n_122), .ZN(p_1[59]));
   OAI21_X1 i_182 (.A(n_123), .B1(n_171), .B2(n_145), .ZN(n_122));
   NAND3_X1 i_183 (.A1(n_146), .A2(n_124), .A3(n_126), .ZN(n_123));
   NOR2_X1 i_184 (.A1(n_173), .A2(n_149), .ZN(n_124));
   INV_X1 i_185 (.A(n_126), .ZN(n_125));
   OAI22_X1 i_186 (.A1(p_0[56]), .A2(aux[56]), .B1(n_150), .B2(n_128), .ZN(n_126));
   OAI21_X1 i_187 (.A(n_151), .B1(p_0[56]), .B2(aux[56]), .ZN(n_127));
   OAI21_X1 i_188 (.A(n_153), .B1(n_175), .B2(n_160), .ZN(n_128));
   AOI21_X1 i_189 (.A(n_174), .B1(p_0[59]), .B2(aux[59]), .ZN(n_129));
   XNOR2_X1 i_190 (.A(n_143), .B(n_142), .ZN(p_1[60]));
   AOI22_X1 i_191 (.A1(n_140), .A2(n_136), .B1(n_141), .B2(n_135), .ZN(p_1[61]));
   XOR2_X1 i_192 (.A(n_131), .B(n_130), .Z(p_1[62]));
   AOI22_X1 i_193 (.A1(p_0[61]), .A2(aux[61]), .B1(n_141), .B2(n_137), .ZN(n_130));
   OAI21_X1 i_194 (.A(n_139), .B1(p_0[62]), .B2(aux[62]), .ZN(n_131));
   XOR2_X1 i_195 (.A(n_133), .B(n_132), .Z(p_1[63]));
   XNOR2_X1 i_196 (.A(p_0[63]), .B(aux[63]), .ZN(n_132));
   OAI221_X1 i_197 (.A(n_134), .B1(p_0[62]), .B2(aux[62]), .C1(n_138), .C2(n_137), 
      .ZN(n_133));
   NAND3_X1 i_198 (.A1(n_139), .A2(n_135), .A3(n_140), .ZN(n_134));
   INV_X1 i_199 (.A(n_136), .ZN(n_135));
   OAI21_X1 i_200 (.A(n_137), .B1(n_379), .B2(n_375), .ZN(n_136));
   NAND2_X1 i_201 (.A1(n_379), .A2(n_375), .ZN(n_137));
   INV_X1 i_202 (.A(n_139), .ZN(n_138));
   NAND2_X1 i_203 (.A1(p_0[62]), .A2(aux[62]), .ZN(n_139));
   INV_X1 i_204 (.A(n_141), .ZN(n_140));
   AOI21_X1 i_205 (.A(n_371), .B1(n_143), .B2(n_142), .ZN(n_141));
   AOI21_X1 i_206 (.A(n_371), .B1(p_0[60]), .B2(aux[60]), .ZN(n_142));
   NOR4_X1 i_207 (.A1(n_147), .A2(n_144), .A3(n_152), .A4(n_159), .ZN(n_143));
   OAI22_X1 i_208 (.A1(n_378), .A2(n_374), .B1(n_174), .B2(n_146), .ZN(n_144));
   INV_X1 i_209 (.A(n_146), .ZN(n_145));
   NAND2_X1 i_210 (.A1(p_0[58]), .A2(aux[58]), .ZN(n_146));
   INV_X1 i_211 (.A(n_148), .ZN(n_147));
   OAI21_X1 i_212 (.A(n_170), .B1(n_150), .B2(n_149), .ZN(n_148));
   AND2_X1 i_213 (.A1(p_0[57]), .A2(aux[57]), .ZN(n_149));
   INV_X1 i_214 (.A(n_151), .ZN(n_150));
   NAND2_X1 i_215 (.A1(p_0[56]), .A2(aux[56]), .ZN(n_151));
   NOR2_X1 i_216 (.A1(n_169), .A2(n_153), .ZN(n_152));
   AOI221_X1 i_217 (.A(n_155), .B1(p_0[55]), .B2(aux[55]), .C1(n_167), .C2(n_154), 
      .ZN(n_153));
   AND2_X1 i_218 (.A1(p_0[54]), .A2(aux[54]), .ZN(n_154));
   AOI21_X1 i_219 (.A(n_162), .B1(n_158), .B2(n_157), .ZN(n_155));
   INV_X1 i_220 (.A(n_157), .ZN(n_156));
   NAND2_X1 i_221 (.A1(p_0[53]), .A2(aux[53]), .ZN(n_157));
   NAND2_X1 i_222 (.A1(p_0[52]), .A2(aux[52]), .ZN(n_158));
   NOR3_X1 i_223 (.A1(n_169), .A2(n_160), .A3(n_175), .ZN(n_159));
   OR2_X1 i_224 (.A1(n_162), .A2(n_161), .ZN(n_160));
   NOR2_X1 i_225 (.A1(p_0[52]), .A2(aux[52]), .ZN(n_161));
   NAND3_X1 i_226 (.A1(n_167), .A2(n_163), .A3(n_165), .ZN(n_162));
   INV_X1 i_227 (.A(n_164), .ZN(n_163));
   NOR2_X1 i_228 (.A1(p_0[54]), .A2(aux[54]), .ZN(n_164));
   INV_X1 i_229 (.A(n_166), .ZN(n_165));
   NOR2_X1 i_230 (.A1(p_0[53]), .A2(aux[53]), .ZN(n_166));
   INV_X1 i_231 (.A(n_168), .ZN(n_167));
   NOR2_X1 i_232 (.A1(p_0[55]), .A2(aux[55]), .ZN(n_168));
   OAI21_X1 i_233 (.A(n_170), .B1(p_0[56]), .B2(aux[56]), .ZN(n_169));
   NOR3_X1 i_234 (.A1(n_174), .A2(n_172), .A3(n_173), .ZN(n_170));
   NOR2_X1 i_235 (.A1(n_173), .A2(n_172), .ZN(n_171));
   NOR2_X1 i_236 (.A1(p_0[58]), .A2(aux[58]), .ZN(n_172));
   NOR2_X1 i_237 (.A1(p_0[57]), .A2(aux[57]), .ZN(n_173));
   NOR2_X1 i_238 (.A1(p_0[59]), .A2(aux[59]), .ZN(n_174));
   NOR4_X1 i_239 (.A1(n_179), .A2(n_176), .A3(n_180), .A4(n_183), .ZN(n_175));
   NOR2_X1 i_240 (.A1(n_188), .A2(n_178), .ZN(n_176));
   INV_X1 i_241 (.A(n_178), .ZN(n_177));
   NAND2_X1 i_242 (.A1(p_0[50]), .A2(aux[50]), .ZN(n_178));
   AND2_X1 i_243 (.A1(p_0[51]), .A2(aux[51]), .ZN(n_179));
   AOI21_X1 i_244 (.A(n_185), .B1(n_182), .B2(n_181), .ZN(n_180));
   NAND2_X1 i_245 (.A1(p_0[49]), .A2(aux[49]), .ZN(n_181));
   NAND2_X1 i_246 (.A1(p_0[48]), .A2(aux[48]), .ZN(n_182));
   NOR3_X1 i_247 (.A1(n_185), .A2(n_184), .A3(n_189), .ZN(n_183));
   NOR2_X1 i_248 (.A1(p_0[48]), .A2(aux[48]), .ZN(n_184));
   OR3_X1 i_249 (.A1(n_188), .A2(n_186), .A3(n_187), .ZN(n_185));
   NOR2_X1 i_250 (.A1(p_0[50]), .A2(aux[50]), .ZN(n_186));
   NOR2_X1 i_251 (.A1(p_0[49]), .A2(aux[49]), .ZN(n_187));
   NOR2_X1 i_252 (.A1(p_0[51]), .A2(aux[51]), .ZN(n_188));
   NOR3_X1 i_253 (.A1(n_211), .A2(n_190), .A3(n_218), .ZN(n_189));
   OAI221_X1 i_254 (.A(n_197), .B1(n_239), .B2(n_191), .C1(n_229), .C2(n_205), 
      .ZN(n_190));
   AOI221_X1 i_255 (.A(n_193), .B1(p_0[43]), .B2(aux[43]), .C1(n_237), .C2(n_192), 
      .ZN(n_191));
   AND2_X1 i_256 (.A1(p_0[42]), .A2(aux[42]), .ZN(n_192));
   AOI21_X1 i_257 (.A(n_232), .B1(n_196), .B2(n_195), .ZN(n_193));
   INV_X1 i_258 (.A(n_195), .ZN(n_194));
   NAND2_X1 i_259 (.A1(p_0[41]), .A2(aux[41]), .ZN(n_195));
   NAND2_X1 i_260 (.A1(p_0[40]), .A2(aux[40]), .ZN(n_196));
   AOI21_X1 i_261 (.A(n_198), .B1(p_0[47]), .B2(aux[47]), .ZN(n_197));
   OAI21_X1 i_262 (.A(n_201), .B1(n_244), .B2(n_200), .ZN(n_198));
   INV_X1 i_263 (.A(n_200), .ZN(n_199));
   NAND2_X1 i_264 (.A1(p_0[46]), .A2(aux[46]), .ZN(n_200));
   OAI21_X1 i_265 (.A(n_240), .B1(n_203), .B2(n_202), .ZN(n_201));
   AND2_X1 i_266 (.A1(p_0[45]), .A2(aux[45]), .ZN(n_202));
   INV_X1 i_267 (.A(n_204), .ZN(n_203));
   NAND2_X1 i_268 (.A1(p_0[44]), .A2(aux[44]), .ZN(n_204));
   AOI221_X1 i_269 (.A(n_207), .B1(p_0[39]), .B2(aux[39]), .C1(n_251), .C2(n_206), 
      .ZN(n_205));
   AND2_X1 i_270 (.A1(p_0[38]), .A2(aux[38]), .ZN(n_206));
   AOI21_X1 i_271 (.A(n_246), .B1(n_210), .B2(n_209), .ZN(n_207));
   INV_X1 i_272 (.A(n_209), .ZN(n_208));
   NAND2_X1 i_273 (.A1(p_0[37]), .A2(aux[37]), .ZN(n_209));
   NAND2_X1 i_274 (.A1(p_0[36]), .A2(aux[36]), .ZN(n_210));
   NOR2_X1 i_275 (.A1(n_228), .A2(n_212), .ZN(n_211));
   AOI221_X1 i_276 (.A(n_214), .B1(p_0[35]), .B2(aux[35]), .C1(n_226), .C2(n_213), 
      .ZN(n_212));
   AND2_X1 i_277 (.A1(p_0[34]), .A2(aux[34]), .ZN(n_213));
   AOI21_X1 i_278 (.A(n_221), .B1(n_217), .B2(n_216), .ZN(n_214));
   INV_X1 i_279 (.A(n_216), .ZN(n_215));
   NAND2_X1 i_280 (.A1(p_0[33]), .A2(aux[33]), .ZN(n_216));
   NAND2_X1 i_281 (.A1(p_0[32]), .A2(aux[32]), .ZN(n_217));
   NOR3_X1 i_282 (.A1(n_228), .A2(n_219), .A3(n_254), .ZN(n_218));
   OR2_X1 i_283 (.A1(n_221), .A2(n_220), .ZN(n_219));
   NOR2_X1 i_284 (.A1(p_0[32]), .A2(aux[32]), .ZN(n_220));
   NAND3_X1 i_285 (.A1(n_226), .A2(n_222), .A3(n_224), .ZN(n_221));
   INV_X1 i_286 (.A(n_223), .ZN(n_222));
   NOR2_X1 i_287 (.A1(p_0[34]), .A2(aux[34]), .ZN(n_223));
   INV_X1 i_288 (.A(n_225), .ZN(n_224));
   NOR2_X1 i_289 (.A1(p_0[33]), .A2(aux[33]), .ZN(n_225));
   INV_X1 i_290 (.A(n_227), .ZN(n_226));
   NOR2_X1 i_291 (.A1(p_0[35]), .A2(aux[35]), .ZN(n_227));
   OR2_X1 i_292 (.A1(n_245), .A2(n_229), .ZN(n_228));
   OR2_X1 i_293 (.A1(n_239), .A2(n_230), .ZN(n_229));
   OR2_X1 i_294 (.A1(n_232), .A2(n_231), .ZN(n_230));
   NOR2_X1 i_295 (.A1(p_0[40]), .A2(aux[40]), .ZN(n_231));
   NAND3_X1 i_296 (.A1(n_237), .A2(n_233), .A3(n_235), .ZN(n_232));
   INV_X1 i_297 (.A(n_234), .ZN(n_233));
   NOR2_X1 i_298 (.A1(p_0[42]), .A2(aux[42]), .ZN(n_234));
   INV_X1 i_299 (.A(n_236), .ZN(n_235));
   NOR2_X1 i_300 (.A1(p_0[41]), .A2(aux[41]), .ZN(n_236));
   INV_X1 i_301 (.A(n_238), .ZN(n_237));
   NOR2_X1 i_302 (.A1(p_0[43]), .A2(aux[43]), .ZN(n_238));
   OAI21_X1 i_303 (.A(n_240), .B1(p_0[44]), .B2(aux[44]), .ZN(n_239));
   NOR3_X1 i_304 (.A1(n_244), .A2(n_242), .A3(n_243), .ZN(n_240));
   NOR2_X1 i_305 (.A1(n_243), .A2(n_242), .ZN(n_241));
   NOR2_X1 i_306 (.A1(p_0[46]), .A2(aux[46]), .ZN(n_242));
   NOR2_X1 i_307 (.A1(p_0[45]), .A2(aux[45]), .ZN(n_243));
   NOR2_X1 i_308 (.A1(p_0[47]), .A2(aux[47]), .ZN(n_244));
   OR2_X1 i_309 (.A1(n_253), .A2(n_246), .ZN(n_245));
   NAND3_X1 i_310 (.A1(n_251), .A2(n_247), .A3(n_249), .ZN(n_246));
   INV_X1 i_311 (.A(n_248), .ZN(n_247));
   NOR2_X1 i_312 (.A1(p_0[38]), .A2(aux[38]), .ZN(n_248));
   INV_X1 i_313 (.A(n_250), .ZN(n_249));
   NOR2_X1 i_314 (.A1(p_0[37]), .A2(aux[37]), .ZN(n_250));
   INV_X1 i_315 (.A(n_252), .ZN(n_251));
   NOR2_X1 i_316 (.A1(p_0[39]), .A2(aux[39]), .ZN(n_252));
   NOR2_X1 i_317 (.A1(p_0[36]), .A2(aux[36]), .ZN(n_253));
   NOR3_X1 i_318 (.A1(n_262), .A2(n_255), .A3(n_280), .ZN(n_254));
   OAI222_X1 i_319 (.A1(n_290), .A2(n_274), .B1(n_291), .B2(n_256), .C1(n_301), 
      .C2(n_268), .ZN(n_255));
   AOI221_X1 i_320 (.A(n_258), .B1(p_0[23]), .B2(aux[23]), .C1(n_316), .C2(n_257), 
      .ZN(n_256));
   AND2_X1 i_321 (.A1(p_0[22]), .A2(aux[22]), .ZN(n_257));
   AOI21_X1 i_322 (.A(n_311), .B1(n_261), .B2(n_260), .ZN(n_258));
   INV_X1 i_323 (.A(n_260), .ZN(n_259));
   NAND2_X1 i_324 (.A1(p_0[21]), .A2(aux[21]), .ZN(n_260));
   NAND2_X1 i_325 (.A1(p_0[20]), .A2(aux[20]), .ZN(n_261));
   OAI222_X1 i_326 (.A1(n_303), .A2(n_265), .B1(n_309), .B2(n_264), .C1(n_377), 
      .C2(n_373), .ZN(n_262));
   INV_X1 i_327 (.A(n_264), .ZN(n_263));
   NAND2_X1 i_328 (.A1(p_0[30]), .A2(aux[30]), .ZN(n_264));
   AOI21_X1 i_329 (.A(n_266), .B1(p_0[28]), .B2(aux[28]), .ZN(n_265));
   AND2_X1 i_330 (.A1(p_0[29]), .A2(aux[29]), .ZN(n_266));
   NAND2_X1 i_331 (.A1(p_0[28]), .A2(aux[28]), .ZN(n_267));
   AOI221_X1 i_332 (.A(n_270), .B1(p_0[27]), .B2(aux[27]), .C1(n_299), .C2(n_269), 
      .ZN(n_268));
   AND2_X1 i_333 (.A1(p_0[26]), .A2(aux[26]), .ZN(n_269));
   AOI21_X1 i_334 (.A(n_294), .B1(n_273), .B2(n_272), .ZN(n_270));
   INV_X1 i_335 (.A(n_272), .ZN(n_271));
   NAND2_X1 i_336 (.A1(p_0[25]), .A2(aux[25]), .ZN(n_272));
   NAND2_X1 i_337 (.A1(p_0[24]), .A2(aux[24]), .ZN(n_273));
   AOI221_X1 i_338 (.A(n_276), .B1(p_0[19]), .B2(aux[19]), .C1(n_288), .C2(n_275), 
      .ZN(n_274));
   AND2_X1 i_339 (.A1(p_0[18]), .A2(aux[18]), .ZN(n_275));
   AOI21_X1 i_340 (.A(n_283), .B1(n_279), .B2(n_278), .ZN(n_276));
   INV_X1 i_341 (.A(n_278), .ZN(n_277));
   NAND2_X1 i_342 (.A1(p_0[17]), .A2(aux[17]), .ZN(n_278));
   NAND2_X1 i_343 (.A1(p_0[16]), .A2(aux[16]), .ZN(n_279));
   NOR3_X1 i_344 (.A1(n_290), .A2(n_281), .A3(n_319), .ZN(n_280));
   OR2_X1 i_345 (.A1(n_283), .A2(n_282), .ZN(n_281));
   NOR2_X1 i_346 (.A1(p_0[16]), .A2(aux[16]), .ZN(n_282));
   NAND3_X1 i_347 (.A1(n_288), .A2(n_284), .A3(n_286), .ZN(n_283));
   INV_X1 i_348 (.A(n_285), .ZN(n_284));
   NOR2_X1 i_349 (.A1(p_0[18]), .A2(aux[18]), .ZN(n_285));
   INV_X1 i_350 (.A(n_287), .ZN(n_286));
   NOR2_X1 i_351 (.A1(p_0[17]), .A2(aux[17]), .ZN(n_287));
   INV_X1 i_352 (.A(n_289), .ZN(n_288));
   NOR2_X1 i_353 (.A1(p_0[19]), .A2(aux[19]), .ZN(n_289));
   OR2_X1 i_354 (.A1(n_310), .A2(n_291), .ZN(n_290));
   OR2_X1 i_355 (.A1(n_301), .A2(n_292), .ZN(n_291));
   OR2_X1 i_356 (.A1(n_294), .A2(n_293), .ZN(n_292));
   NOR2_X1 i_357 (.A1(p_0[24]), .A2(aux[24]), .ZN(n_293));
   NAND3_X1 i_358 (.A1(n_299), .A2(n_295), .A3(n_297), .ZN(n_294));
   INV_X1 i_359 (.A(n_296), .ZN(n_295));
   NOR2_X1 i_360 (.A1(p_0[26]), .A2(aux[26]), .ZN(n_296));
   INV_X1 i_361 (.A(n_298), .ZN(n_297));
   NOR2_X1 i_362 (.A1(p_0[25]), .A2(aux[25]), .ZN(n_298));
   INV_X1 i_363 (.A(n_300), .ZN(n_299));
   NOR2_X1 i_364 (.A1(p_0[27]), .A2(aux[27]), .ZN(n_300));
   OR2_X1 i_365 (.A1(n_303), .A2(n_302), .ZN(n_301));
   NOR2_X1 i_366 (.A1(p_0[28]), .A2(aux[28]), .ZN(n_302));
   NAND3_X1 i_367 (.A1(n_308), .A2(n_304), .A3(n_306), .ZN(n_303));
   INV_X1 i_368 (.A(n_305), .ZN(n_304));
   NOR2_X1 i_369 (.A1(p_0[30]), .A2(aux[30]), .ZN(n_305));
   INV_X1 i_370 (.A(n_307), .ZN(n_306));
   NOR2_X1 i_371 (.A1(p_0[29]), .A2(aux[29]), .ZN(n_307));
   INV_X1 i_372 (.A(n_309), .ZN(n_308));
   NOR2_X1 i_373 (.A1(p_0[31]), .A2(aux[31]), .ZN(n_309));
   OR2_X1 i_374 (.A1(n_318), .A2(n_311), .ZN(n_310));
   NAND3_X1 i_375 (.A1(n_316), .A2(n_312), .A3(n_314), .ZN(n_311));
   INV_X1 i_376 (.A(n_313), .ZN(n_312));
   NOR2_X1 i_377 (.A1(p_0[22]), .A2(aux[22]), .ZN(n_313));
   INV_X1 i_378 (.A(n_315), .ZN(n_314));
   NOR2_X1 i_379 (.A1(p_0[21]), .A2(aux[21]), .ZN(n_315));
   INV_X1 i_380 (.A(n_317), .ZN(n_316));
   NOR2_X1 i_381 (.A1(p_0[23]), .A2(aux[23]), .ZN(n_317));
   NOR2_X1 i_382 (.A1(p_0[20]), .A2(aux[20]), .ZN(n_318));
   NOR4_X1 i_383 (.A1(n_323), .A2(n_320), .A3(n_324), .A4(n_327), .ZN(n_319));
   NOR2_X1 i_384 (.A1(n_332), .A2(n_322), .ZN(n_320));
   INV_X1 i_385 (.A(n_322), .ZN(n_321));
   NAND2_X1 i_386 (.A1(p_0[14]), .A2(aux[14]), .ZN(n_322));
   AND2_X1 i_387 (.A1(p_0[15]), .A2(aux[15]), .ZN(n_323));
   AOI21_X1 i_388 (.A(n_329), .B1(n_326), .B2(n_325), .ZN(n_324));
   NAND2_X1 i_389 (.A1(p_0[13]), .A2(aux[13]), .ZN(n_325));
   NAND2_X1 i_390 (.A1(p_0[12]), .A2(aux[12]), .ZN(n_326));
   NOR3_X1 i_391 (.A1(n_329), .A2(n_328), .A3(n_333), .ZN(n_327));
   NOR2_X1 i_392 (.A1(p_0[12]), .A2(aux[12]), .ZN(n_328));
   OR3_X1 i_393 (.A1(n_332), .A2(n_330), .A3(n_331), .ZN(n_329));
   NOR2_X1 i_394 (.A1(p_0[14]), .A2(aux[14]), .ZN(n_330));
   NOR2_X1 i_395 (.A1(p_0[13]), .A2(aux[13]), .ZN(n_331));
   NOR2_X1 i_396 (.A1(p_0[15]), .A2(aux[15]), .ZN(n_332));
   NOR4_X1 i_397 (.A1(n_337), .A2(n_334), .A3(n_338), .A4(n_341), .ZN(n_333));
   NOR2_X1 i_398 (.A1(n_346), .A2(n_336), .ZN(n_334));
   INV_X1 i_399 (.A(n_336), .ZN(n_335));
   NAND2_X1 i_400 (.A1(p_0[10]), .A2(aux[10]), .ZN(n_336));
   AND2_X1 i_401 (.A1(p_0[11]), .A2(aux[11]), .ZN(n_337));
   AOI21_X1 i_402 (.A(n_343), .B1(n_340), .B2(n_339), .ZN(n_338));
   NAND2_X1 i_403 (.A1(p_0[9]), .A2(aux[9]), .ZN(n_339));
   NAND2_X1 i_404 (.A1(p_0[8]), .A2(aux[8]), .ZN(n_340));
   NOR3_X1 i_405 (.A1(n_343), .A2(n_342), .A3(n_347), .ZN(n_341));
   NOR2_X1 i_406 (.A1(p_0[8]), .A2(aux[8]), .ZN(n_342));
   OR3_X1 i_407 (.A1(n_346), .A2(n_344), .A3(n_345), .ZN(n_343));
   NOR2_X1 i_408 (.A1(p_0[10]), .A2(aux[10]), .ZN(n_344));
   NOR2_X1 i_409 (.A1(p_0[9]), .A2(aux[9]), .ZN(n_345));
   NOR2_X1 i_410 (.A1(p_0[11]), .A2(aux[11]), .ZN(n_346));
   NOR4_X1 i_411 (.A1(n_351), .A2(n_348), .A3(n_352), .A4(n_355), .ZN(n_347));
   NOR2_X1 i_412 (.A1(n_360), .A2(n_350), .ZN(n_348));
   INV_X1 i_413 (.A(n_350), .ZN(n_349));
   NAND2_X1 i_414 (.A1(p_0[6]), .A2(aux[6]), .ZN(n_350));
   AND2_X1 i_415 (.A1(p_0[7]), .A2(aux[7]), .ZN(n_351));
   AOI21_X1 i_416 (.A(n_357), .B1(n_354), .B2(n_353), .ZN(n_352));
   NAND2_X1 i_417 (.A1(p_0[5]), .A2(aux[5]), .ZN(n_353));
   NAND2_X1 i_418 (.A1(p_0[4]), .A2(aux[4]), .ZN(n_354));
   NOR3_X1 i_419 (.A1(n_357), .A2(n_356), .A3(n_361), .ZN(n_355));
   NOR2_X1 i_420 (.A1(p_0[4]), .A2(aux[4]), .ZN(n_356));
   OR3_X1 i_421 (.A1(n_360), .A2(n_358), .A3(n_359), .ZN(n_357));
   NOR2_X1 i_422 (.A1(p_0[6]), .A2(aux[6]), .ZN(n_358));
   NOR2_X1 i_423 (.A1(p_0[5]), .A2(aux[5]), .ZN(n_359));
   NOR2_X1 i_424 (.A1(p_0[7]), .A2(aux[7]), .ZN(n_360));
   NAND2_X1 i_425 (.A1(n_370), .A2(n_362), .ZN(n_361));
   OAI21_X1 i_426 (.A(n_363), .B1(n_376), .B2(n_372), .ZN(n_362));
   OAI22_X1 i_427 (.A1(p_0[2]), .A2(aux[2]), .B1(n_368), .B2(n_364), .ZN(n_363));
   AOI21_X1 i_428 (.A(n_367), .B1(n_366), .B2(n_365), .ZN(n_364));
   NAND2_X1 i_429 (.A1(p_0[1]), .A2(aux[1]), .ZN(n_365));
   NAND2_X1 i_430 (.A1(p_0[0]), .A2(aux[0]), .ZN(n_366));
   NOR2_X1 i_431 (.A1(p_0[1]), .A2(aux[1]), .ZN(n_367));
   INV_X1 i_432 (.A(n_369), .ZN(n_368));
   NAND2_X1 i_433 (.A1(p_0[2]), .A2(aux[2]), .ZN(n_369));
   NAND2_X1 i_434 (.A1(n_376), .A2(n_372), .ZN(n_370));
   NOR2_X1 i_435 (.A1(p_0[60]), .A2(aux[60]), .ZN(n_371));
   INV_X1 i_436 (.A(aux[3]), .ZN(n_372));
   INV_X1 i_437 (.A(aux[31]), .ZN(n_373));
   INV_X1 i_438 (.A(aux[59]), .ZN(n_374));
   INV_X1 i_439 (.A(aux[61]), .ZN(n_375));
   INV_X1 i_440 (.A(p_0[3]), .ZN(n_376));
   INV_X1 i_441 (.A(p_0[31]), .ZN(n_377));
   INV_X1 i_442 (.A(p_0[59]), .ZN(n_378));
   INV_X1 i_443 (.A(p_0[61]), .ZN(n_379));
endmodule

module radix4Booth(a, b, clk, reset, en, result, enableOutput);
   input [31:0]a;
   input [31:0]b;
   input clk;
   input reset;
   input en;
   output [63:0]result;
   output enableOutput;

   wire [31:0]firstInputComplement;
   wire n_1_3;
   wire n_1_0;
   wire n_1_4;
   wire n_1_1;
   wire n_1_5;
   wire n_1_2;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_115;
   wire n_1_116;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_123;
   wire n_1_124;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_149;
   wire n_1_150;
   wire n_1_151;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_160;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_169;
   wire n_1_170;
   wire n_1_171;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;
   wire n_1_176;
   wire n_1_177;
   wire n_1_178;
   wire n_1_179;
   wire n_1_180;
   wire n_1_181;
   wire n_1_182;
   wire n_1_183;
   wire n_1_184;
   wire n_1_185;
   wire n_1_186;
   wire n_1_187;
   wire n_1_188;
   wire n_1_189;
   wire n_1_190;
   wire n_1_191;
   wire n_1_192;
   wire n_1_193;
   wire n_1_194;
   wire n_1_195;
   wire n_1_196;
   wire n_1_197;
   wire n_1_198;
   wire n_1_199;
   wire n_1_200;
   wire n_1_201;
   wire n_1_202;
   wire n_1_203;
   wire n_1_204;
   wire n_1_205;
   wire n_1_206;
   wire n_1_207;
   wire n_1_208;
   wire n_1_209;
   wire n_1_210;
   wire n_1_211;
   wire n_1_212;
   wire n_1_213;
   wire n_1_214;
   wire n_1_215;
   wire n_1_216;
   wire n_1_217;
   wire n_1_218;
   wire n_1_219;
   wire n_1_220;
   wire n_1_221;
   wire n_1_222;
   wire n_1_223;
   wire n_1_224;
   wire n_1_225;
   wire n_1_226;
   wire n_1_227;
   wire n_1_228;
   wire n_1_229;
   wire n_1_230;
   wire n_1_231;
   wire n_1_232;
   wire n_1_233;
   wire n_1_234;
   wire n_1_235;
   wire n_1_236;
   wire n_1_237;
   wire n_1_238;
   wire n_1_239;
   wire n_1_240;
   wire n_1_241;
   wire n_1_242;
   wire n_1_243;
   wire n_1_244;
   wire n_1_245;
   wire n_1_246;
   wire n_1_247;
   wire n_1_248;
   wire n_1_249;
   wire n_1_250;
   wire n_1_251;
   wire n_1_252;
   wire n_1_253;
   wire n_1_254;
   wire n_1_255;
   wire n_1_256;
   wire n_1_257;
   wire n_1_258;
   wire n_1_259;
   wire n_1_260;
   wire n_1_261;
   wire n_1_262;
   wire n_1_263;
   wire n_1_264;
   wire n_1_265;
   wire n_1_266;
   wire n_1_267;
   wire n_1_268;
   wire n_1_269;
   wire n_1_270;
   wire n_1_271;
   wire n_1_272;
   wire n_1_273;
   wire n_1_274;
   wire n_1_275;
   wire n_1_276;
   wire n_1_277;
   wire n_1_278;
   wire n_1_279;
   wire n_1_280;
   wire n_1_281;
   wire n_1_282;
   wire n_1_283;
   wire n_1_284;
   wire n_1_285;
   wire n_1_286;
   wire n_1_287;
   wire n_1_288;
   wire n_1_289;
   wire n_1_290;
   wire n_1_291;
   wire n_1_292;
   wire n_1_293;
   wire n_1_294;
   wire n_1_295;
   wire n_1_296;
   wire n_1_297;
   wire n_1_298;
   wire n_1_299;
   wire n_1_300;
   wire n_1_301;
   wire n_1_302;
   wire n_1_303;
   wire n_1_304;
   wire n_1_305;
   wire n_1_306;
   wire n_1_307;
   wire n_1_308;
   wire n_1_309;
   wire n_1_310;
   wire n_1_311;
   wire n_1_312;
   wire n_1_313;
   wire n_1_314;
   wire n_1_315;
   wire n_1_316;
   wire n_1_317;
   wire n_1_318;
   wire n_1_319;
   wire n_1_320;
   wire n_1_321;
   wire n_1_322;
   wire n_1_323;
   wire n_1_324;
   wire n_1_325;
   wire n_1_326;
   wire n_1_327;
   wire n_1_328;
   wire n_1_329;
   wire n_1_330;
   wire n_1_331;
   wire n_1_332;
   wire n_1_333;
   wire n_1_334;
   wire n_1_335;
   wire n_1_336;
   wire n_1_337;
   wire n_1_338;
   wire n_1_339;
   wire n_1_340;
   wire n_1_341;
   wire n_1_342;
   wire n_1_343;
   wire n_1_344;
   wire n_1_345;
   wire n_1_346;
   wire n_1_347;
   wire n_1_348;
   wire n_1_349;
   wire n_1_350;
   wire n_1_351;
   wire n_1_352;
   wire n_1_353;
   wire n_1_354;
   wire n_1_355;
   wire n_1_356;
   wire n_1_357;
   wire n_1_358;
   wire n_1_359;
   wire n_1_360;
   wire n_1_361;
   wire n_1_362;
   wire n_1_363;
   wire n_1_364;
   wire n_1_365;
   wire n_1_366;
   wire n_1_367;
   wire n_1_368;
   wire n_1_369;
   wire n_1_370;
   wire n_1_371;
   wire n_1_372;
   wire n_1_373;
   wire n_1_374;
   wire n_1_375;
   wire n_1_376;
   wire n_1_377;
   wire n_1_378;
   wire n_1_379;
   wire n_1_380;
   wire n_1_381;
   wire n_1_382;
   wire n_1_383;
   wire n_1_384;
   wire n_1_385;
   wire n_1_386;
   wire n_1_387;
   wire n_1_388;
   wire n_1_389;
   wire n_1_390;
   wire n_1_391;
   wire n_1_392;
   wire n_1_393;
   wire n_1_394;
   wire n_1_395;
   wire n_1_396;
   wire n_1_397;
   wire n_1_398;
   wire n_1_399;
   wire n_1_400;
   wire n_1_401;
   wire n_1_402;
   wire n_1_403;
   wire n_1_404;
   wire n_1_405;
   wire n_1_406;
   wire n_1_407;
   wire n_1_408;
   wire n_1_409;
   wire n_1_410;
   wire n_1_411;
   wire n_1_412;
   wire n_1_413;
   wire n_1_414;
   wire n_1_415;
   wire n_1_416;
   wire n_1_417;
   wire n_1_418;
   wire n_1_419;
   wire n_1_420;
   wire n_1_421;
   wire n_1_422;
   wire n_1_423;
   wire n_1_424;
   wire n_1_425;
   wire n_1_426;
   wire n_1_427;
   wire n_1_428;
   wire n_1_429;
   wire n_1_430;
   wire n_1_431;
   wire n_1_432;
   wire n_1_433;
   wire n_1_434;
   wire n_1_435;
   wire n_1_436;
   wire n_1_437;
   wire n_1_438;
   wire n_1_439;
   wire n_1_440;
   wire n_1_441;
   wire n_1_442;
   wire n_1_443;
   wire n_1_444;
   wire n_1_445;
   wire n_1_446;
   wire n_1_447;
   wire n_1_448;
   wire n_1_449;
   wire n_1_450;
   wire n_1_451;
   wire n_1_452;
   wire n_1_453;
   wire n_1_454;
   wire n_1_455;
   wire n_1_456;
   wire n_1_457;
   wire n_1_458;
   wire n_1_459;
   wire n_1_460;
   wire n_1_461;
   wire n_1_462;
   wire n_1_463;
   wire n_1_464;
   wire n_1_465;
   wire n_1_466;
   wire n_1_467;
   wire n_1_468;
   wire n_1_469;
   wire n_1_470;
   wire n_1_471;
   wire n_1_472;
   wire n_1_473;
   wire n_1_474;
   wire n_1_475;
   wire n_1_476;
   wire n_1_477;
   wire n_1_478;
   wire n_1_479;
   wire n_1_480;
   wire n_1_481;
   wire n_1_482;
   wire n_1_483;
   wire n_1_484;
   wire n_1_485;
   wire n_1_486;
   wire n_1_487;
   wire n_1_488;
   wire n_1_489;
   wire n_1_490;
   wire n_1_491;
   wire n_1_492;
   wire n_1_493;
   wire n_1_494;
   wire n_1_495;
   wire n_1_496;
   wire n_1_497;
   wire n_1_498;
   wire n_1_499;
   wire n_1_500;
   wire n_1_501;
   wire n_1_502;
   wire n_1_503;
   wire n_1_504;
   wire n_1_505;
   wire n_1_506;
   wire n_1_507;
   wire n_1_508;
   wire n_1_509;
   wire n_1_510;
   wire n_1_511;
   wire n_1_512;
   wire n_1_513;
   wire n_1_514;
   wire n_1_515;
   wire n_1_516;
   wire n_1_517;
   wire n_1_518;
   wire n_1_519;
   wire n_1_520;
   wire n_1_521;
   wire n_1_522;
   wire n_1_523;
   wire n_1_524;
   wire n_1_525;
   wire n_1_526;
   wire n_1_527;
   wire n_1_528;
   wire n_1_529;
   wire n_1_530;
   wire n_1_531;
   wire n_1_532;
   wire n_1_533;
   wire n_1_534;
   wire n_1_535;
   wire n_1_536;
   wire n_1_537;
   wire n_1_538;
   wire n_1_539;
   wire n_1_540;
   wire n_1_541;
   wire n_1_542;
   wire n_1_543;
   wire n_1_544;
   wire n_1_545;
   wire n_1_546;
   wire n_1_547;
   wire n_1_548;
   wire n_1_549;
   wire n_1_550;
   wire n_1_551;
   wire n_1_552;
   wire n_1_553;
   wire n_1_554;
   wire n_1_555;
   wire n_1_556;
   wire n_1_557;
   wire n_1_558;
   wire n_1_559;
   wire n_1_560;
   wire n_1_561;
   wire n_1_562;
   wire n_1_563;
   wire n_1_564;
   wire n_1_565;
   wire n_1_566;
   wire n_1_567;
   wire n_1_568;
   wire n_1_569;
   wire n_1_570;
   wire n_1_571;
   wire n_1_572;
   wire n_1_573;
   wire n_1_574;
   wire n_1_575;
   wire n_1_576;
   wire n_1_577;
   wire n_1_578;
   wire n_1_579;
   wire n_1_580;
   wire n_1_581;
   wire n_1_582;
   wire n_1_583;
   wire n_1_584;
   wire n_1_585;
   wire n_1_586;
   wire n_1_587;
   wire n_1_588;
   wire n_1_589;
   wire n_1_590;
   wire n_1_591;
   wire n_1_592;
   wire n_1_593;
   wire n_1_594;
   wire n_1_595;
   wire n_1_596;
   wire n_1_597;
   wire n_1_598;
   wire n_1_599;
   wire n_1_600;
   wire n_1_601;
   wire n_1_602;
   wire n_1_603;
   wire n_1_604;
   wire n_1_605;
   wire n_1_606;
   wire n_1_607;
   wire n_1_608;
   wire n_1_609;
   wire n_1_610;
   wire n_1_611;
   wire n_1_612;
   wire n_1_613;
   wire n_1_614;
   wire n_1_615;
   wire n_1_616;
   wire n_1_617;
   wire n_1_618;
   wire n_1_619;
   wire n_1_620;
   wire n_1_621;
   wire n_1_622;
   wire n_1_623;
   wire n_1_624;
   wire n_1_625;
   wire n_1_626;
   wire n_1_627;
   wire n_1_628;
   wire n_1_629;
   wire n_1_630;
   wire n_1_631;
   wire n_1_632;
   wire n_1_633;
   wire n_1_634;
   wire n_1_635;
   wire n_1_636;
   wire n_1_637;
   wire n_1_638;
   wire n_1_639;
   wire n_1_640;
   wire n_1_641;
   wire n_1_642;
   wire n_1_643;
   wire n_1_644;
   wire n_1_645;
   wire n_1_646;
   wire n_1_647;
   wire n_1_648;
   wire n_1_649;
   wire n_1_650;
   wire n_1_651;
   wire n_1_652;
   wire n_1_653;
   wire n_1_654;
   wire n_1_655;
   wire n_1_656;
   wire n_1_657;
   wire n_1_658;
   wire n_1_659;
   wire n_1_660;
   wire n_1_661;
   wire n_1_662;
   wire n_1_663;
   wire n_1_664;
   wire n_1_665;
   wire n_1_666;
   wire n_1_667;
   wire n_1_668;
   wire n_1_669;
   wire n_1_670;
   wire n_1_671;
   wire n_1_672;
   wire n_1_673;
   wire n_1_674;
   wire n_1_675;
   wire n_1_676;
   wire n_1_677;
   wire n_1_678;
   wire n_1_679;
   wire n_1_680;
   wire n_1_681;
   wire n_1_682;
   wire n_1_683;
   wire n_1_684;
   wire n_1_685;
   wire n_1_686;
   wire n_1_687;
   wire n_1_688;
   wire n_1_689;
   wire n_1_690;
   wire n_1_691;
   wire n_1_692;
   wire n_1_693;
   wire n_1_694;
   wire n_1_695;
   wire n_1_696;
   wire n_1_697;
   wire n_1_698;
   wire n_1_699;
   wire n_1_700;
   wire n_1_701;
   wire n_1_702;
   wire n_1_703;
   wire n_1_704;
   wire n_1_705;
   wire n_1_706;
   wire n_1_707;
   wire n_1_708;
   wire n_1_709;
   wire n_1_710;
   wire n_1_711;
   wire n_1_712;
   wire n_1_713;
   wire n_1_714;
   wire n_1_715;
   wire n_1_716;
   wire n_1_717;
   wire n_1_718;
   wire n_1_719;
   wire n_1_720;
   wire n_1_721;
   wire n_1_722;
   wire n_1_723;
   wire n_1_724;
   wire n_1_725;
   wire n_1_726;
   wire n_1_727;
   wire n_1_728;
   wire n_1_729;
   wire n_1_730;
   wire n_1_731;
   wire n_1_732;
   wire n_1_733;
   wire n_1_734;
   wire n_1_735;
   wire n_1_736;
   wire n_1_737;
   wire n_1_738;
   wire n_1_739;
   wire n_1_740;
   wire n_1_741;
   wire n_1_742;
   wire n_1_743;
   wire n_1_744;
   wire n_1_745;
   wire n_1_746;
   wire n_1_747;
   wire n_1_748;
   wire n_1_749;
   wire n_1_750;
   wire n_1_751;
   wire n_1_752;
   wire n_1_753;
   wire n_1_754;
   wire n_1_755;
   wire n_1_756;
   wire n_1_757;
   wire n_1_758;
   wire n_1_759;
   wire n_1_760;
   wire n_1_761;
   wire n_1_762;
   wire n_1_763;
   wire n_1_764;
   wire n_1_765;
   wire n_1_766;
   wire n_1_767;
   wire n_1_768;
   wire n_1_769;
   wire n_1_770;
   wire n_1_771;
   wire n_1_772;
   wire n_1_773;
   wire n_1_774;
   wire n_1_775;
   wire n_1_776;
   wire n_1_777;
   wire n_1_778;
   wire n_1_779;
   wire n_1_780;
   wire n_1_781;
   wire n_1_782;
   wire n_1_783;
   wire n_1_784;
   wire n_1_785;
   wire n_1_786;
   wire n_1_787;
   wire n_1_788;
   wire n_1_789;
   wire n_1_790;
   wire n_1_791;
   wire n_1_792;
   wire n_1_793;
   wire n_1_794;
   wire n_1_795;
   wire n_1_796;
   wire n_1_797;
   wire n_1_798;
   wire n_1_799;
   wire n_1_800;
   wire n_1_801;
   wire n_1_802;
   wire n_1_803;
   wire n_1_804;
   wire n_1_805;
   wire n_1_806;
   wire n_1_807;
   wire n_1_808;
   wire n_1_809;
   wire n_1_810;
   wire n_1_811;
   wire n_1_812;
   wire n_1_813;
   wire n_1_814;
   wire n_1_815;
   wire n_1_816;
   wire n_1_817;
   wire n_1_818;
   wire n_1_819;
   wire n_1_820;
   wire n_1_821;
   wire n_1_822;
   wire n_1_823;
   wire n_1_824;
   wire n_1_825;
   wire n_1_826;
   wire n_1_827;
   wire n_1_828;
   wire n_1_829;
   wire n_1_830;
   wire n_1_831;
   wire n_1_832;
   wire n_1_833;
   wire n_1_834;
   wire n_1_835;
   wire n_1_836;
   wire n_1_837;
   wire n_1_838;
   wire n_1_839;
   wire n_1_840;
   wire n_1_841;
   wire n_1_842;
   wire n_1_843;
   wire n_1_844;
   wire n_1_845;
   wire n_1_846;
   wire n_1_847;
   wire n_1_848;
   wire n_1_849;
   wire n_1_850;
   wire n_1_851;
   wire n_1_852;
   wire n_1_853;
   wire n_1_854;
   wire n_1_855;
   wire n_1_856;
   wire n_1_857;
   wire n_1_858;
   wire n_1_859;
   wire n_1_860;
   wire n_1_861;
   wire n_1_862;
   wire n_1_863;
   wire n_1_864;
   wire n_1_865;
   wire n_1_866;
   wire n_1_867;
   wire n_1_868;
   wire n_1_869;
   wire n_1_870;
   wire n_1_871;
   wire n_1_872;
   wire n_1_873;
   wire n_1_874;
   wire n_1_875;
   wire n_1_876;
   wire n_1_877;
   wire n_1_878;
   wire n_1_879;
   wire n_1_880;
   wire n_1_881;
   wire n_1_882;
   wire n_1_883;
   wire n_1_884;
   wire n_1_885;
   wire n_1_886;
   wire n_1_887;
   wire n_1_888;
   wire n_1_889;
   wire n_1_890;
   wire n_1_891;
   wire n_1_892;
   wire n_1_893;
   wire n_1_894;
   wire n_1_895;
   wire n_1_896;
   wire n_1_897;
   wire n_1_898;
   wire n_1_899;
   wire n_1_900;
   wire n_1_901;
   wire n_1_902;
   wire n_1_903;
   wire n_1_904;
   wire n_1_905;
   wire n_1_906;
   wire n_1_907;
   wire n_1_908;
   wire n_1_909;
   wire n_1_910;
   wire n_1_911;
   wire n_1_912;
   wire n_1_913;
   wire n_1_914;
   wire n_1_915;
   wire n_1_916;
   wire n_1_917;
   wire n_1_918;
   wire n_1_919;
   wire n_1_920;
   wire n_1_921;
   wire n_1_922;
   wire n_1_923;
   wire n_1_924;
   wire n_1_925;
   wire n_1_926;
   wire n_1_927;
   wire n_1_928;
   wire n_1_929;
   wire n_1_930;
   wire n_1_931;
   wire n_1_932;
   wire n_1_933;
   wire n_1_934;
   wire n_1_935;
   wire n_1_936;
   wire n_1_937;
   wire n_1_938;
   wire [4:0]counter;
   wire resetReg;
   wire [63:0]aux;

   datapath i_0 (.firstInputComplement({firstInputComplement[31], 
      firstInputComplement[30], firstInputComplement[29], 
      firstInputComplement[28], firstInputComplement[27], 
      firstInputComplement[26], firstInputComplement[25], 
      firstInputComplement[24], firstInputComplement[23], 
      firstInputComplement[22], firstInputComplement[21], 
      firstInputComplement[20], firstInputComplement[19], 
      firstInputComplement[18], firstInputComplement[17], 
      firstInputComplement[16], firstInputComplement[15], 
      firstInputComplement[14], firstInputComplement[13], 
      firstInputComplement[12], firstInputComplement[11], 
      firstInputComplement[10], firstInputComplement[9], firstInputComplement[8], 
      firstInputComplement[7], firstInputComplement[6], firstInputComplement[5], 
      firstInputComplement[4], firstInputComplement[3], firstInputComplement[2], 
      firstInputComplement[1], uc_0}), .a(a));
   DFF_X1 enableOutput_reg (.D(n_268), .CK(clk), .Q(enableOutput), .QN());
   datapath__0_74 i_41 (.p_0({n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
      n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, n_249, n_248, 
      n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, n_238, 
      n_237, n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, n_228, 
      n_227, n_226, n_225, n_224, n_223, n_222, n_221, n_220, n_219, n_218, 
      n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, 
      n_207, n_206, n_205, n_204, n_203, n_202, n_201}), .aux(aux), .p_1({n_66, 
      n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
      n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
      n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
      n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, 
      n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
      n_4, n_3}));
   HA_X1 i_1_0 (.A(counter[1]), .B(counter[0]), .CO(n_1_0), .S(n_1_3));
   HA_X1 i_1_1 (.A(counter[2]), .B(n_1_0), .CO(n_1_1), .S(n_1_4));
   HA_X1 i_1_2 (.A(counter[3]), .B(n_1_1), .CO(n_1_2), .S(n_1_5));
   AND2_X1 i_1_3 (.A1(en), .A2(reset), .ZN(n_67));
   NOR2_X1 i_1_4 (.A1(n_1_795), .A2(n_267), .ZN(n_68));
   NOR2_X1 i_1_5 (.A1(n_1_796), .A2(n_267), .ZN(n_69));
   NOR2_X1 i_1_6 (.A1(n_1_797), .A2(n_267), .ZN(n_70));
   NOR2_X1 i_1_7 (.A1(n_1_798), .A2(n_267), .ZN(n_71));
   NOR2_X1 i_1_8 (.A1(n_1_799), .A2(n_267), .ZN(n_72));
   NOR2_X1 i_1_9 (.A1(n_1_800), .A2(n_267), .ZN(n_73));
   NOR2_X1 i_1_10 (.A1(n_1_801), .A2(n_267), .ZN(n_74));
   NOR2_X1 i_1_11 (.A1(n_1_802), .A2(n_267), .ZN(n_75));
   NOR2_X1 i_1_12 (.A1(n_1_803), .A2(n_267), .ZN(n_76));
   NOR2_X1 i_1_13 (.A1(n_1_804), .A2(n_267), .ZN(n_77));
   NOR2_X1 i_1_14 (.A1(n_1_805), .A2(n_267), .ZN(n_78));
   NOR2_X1 i_1_15 (.A1(n_1_806), .A2(n_267), .ZN(n_79));
   NOR2_X1 i_1_16 (.A1(n_1_807), .A2(n_267), .ZN(n_80));
   NOR2_X1 i_1_17 (.A1(n_1_808), .A2(n_267), .ZN(n_81));
   NOR2_X1 i_1_18 (.A1(n_1_809), .A2(n_267), .ZN(n_82));
   NOR2_X1 i_1_19 (.A1(n_1_810), .A2(n_267), .ZN(n_83));
   NOR2_X1 i_1_20 (.A1(n_1_811), .A2(n_267), .ZN(n_84));
   NOR2_X1 i_1_21 (.A1(n_1_812), .A2(n_267), .ZN(n_85));
   NOR2_X1 i_1_22 (.A1(n_1_813), .A2(n_267), .ZN(n_86));
   NOR2_X1 i_1_23 (.A1(n_1_814), .A2(n_267), .ZN(n_87));
   NOR2_X1 i_1_24 (.A1(n_1_815), .A2(n_267), .ZN(n_88));
   NOR2_X1 i_1_25 (.A1(n_1_816), .A2(n_267), .ZN(n_89));
   NOR2_X1 i_1_26 (.A1(n_1_817), .A2(n_267), .ZN(n_90));
   NOR2_X1 i_1_27 (.A1(n_1_818), .A2(n_267), .ZN(n_91));
   NOR2_X1 i_1_28 (.A1(n_1_819), .A2(n_267), .ZN(n_92));
   NOR2_X1 i_1_29 (.A1(n_1_820), .A2(n_267), .ZN(n_93));
   NOR2_X1 i_1_30 (.A1(n_1_821), .A2(n_267), .ZN(n_94));
   NOR2_X1 i_1_31 (.A1(n_1_822), .A2(n_267), .ZN(n_95));
   NOR2_X1 i_1_32 (.A1(n_1_823), .A2(n_267), .ZN(n_96));
   NOR2_X1 i_1_33 (.A1(n_1_824), .A2(n_267), .ZN(n_97));
   NOR2_X1 i_1_34 (.A1(n_1_825), .A2(n_267), .ZN(n_98));
   NOR2_X1 i_1_35 (.A1(n_1_826), .A2(n_267), .ZN(n_99));
   NOR2_X1 i_1_36 (.A1(n_1_827), .A2(n_267), .ZN(n_100));
   NOR2_X1 i_1_37 (.A1(n_1_828), .A2(n_267), .ZN(n_101));
   NOR2_X1 i_1_38 (.A1(n_1_829), .A2(n_267), .ZN(n_102));
   NOR2_X1 i_1_39 (.A1(n_1_830), .A2(n_267), .ZN(n_103));
   NOR2_X1 i_1_40 (.A1(n_1_831), .A2(n_267), .ZN(n_104));
   NOR2_X1 i_1_41 (.A1(n_1_832), .A2(n_267), .ZN(n_105));
   NOR2_X1 i_1_42 (.A1(n_1_833), .A2(n_267), .ZN(n_106));
   NOR2_X1 i_1_43 (.A1(n_1_834), .A2(n_267), .ZN(n_107));
   NOR2_X1 i_1_44 (.A1(n_1_835), .A2(n_267), .ZN(n_108));
   NOR2_X1 i_1_45 (.A1(n_1_836), .A2(n_267), .ZN(n_109));
   NOR2_X1 i_1_46 (.A1(n_1_837), .A2(n_267), .ZN(n_110));
   NOR2_X1 i_1_47 (.A1(n_1_838), .A2(n_267), .ZN(n_111));
   NOR2_X1 i_1_48 (.A1(n_1_839), .A2(n_267), .ZN(n_112));
   NOR2_X1 i_1_49 (.A1(n_1_840), .A2(n_267), .ZN(n_113));
   NOR2_X1 i_1_50 (.A1(n_1_841), .A2(n_267), .ZN(n_114));
   NOR2_X1 i_1_51 (.A1(n_1_842), .A2(n_267), .ZN(n_115));
   NOR2_X1 i_1_52 (.A1(n_1_843), .A2(n_267), .ZN(n_116));
   NOR2_X1 i_1_53 (.A1(n_1_844), .A2(n_267), .ZN(n_117));
   NOR2_X1 i_1_54 (.A1(n_1_845), .A2(n_267), .ZN(n_118));
   NOR2_X1 i_1_55 (.A1(n_1_846), .A2(n_267), .ZN(n_119));
   NOR2_X1 i_1_56 (.A1(n_1_847), .A2(n_267), .ZN(n_120));
   NOR2_X1 i_1_57 (.A1(n_1_848), .A2(n_267), .ZN(n_121));
   NOR2_X1 i_1_58 (.A1(n_1_849), .A2(n_267), .ZN(n_122));
   NOR2_X1 i_1_59 (.A1(n_1_850), .A2(n_267), .ZN(n_123));
   NOR2_X1 i_1_60 (.A1(n_1_851), .A2(n_267), .ZN(n_124));
   NOR2_X1 i_1_61 (.A1(n_1_852), .A2(n_267), .ZN(n_125));
   NOR2_X1 i_1_62 (.A1(n_1_853), .A2(n_267), .ZN(n_126));
   NOR2_X1 i_1_63 (.A1(n_1_854), .A2(n_267), .ZN(n_127));
   NOR2_X1 i_1_64 (.A1(n_1_855), .A2(n_267), .ZN(n_128));
   NOR2_X1 i_1_65 (.A1(n_1_856), .A2(n_267), .ZN(n_129));
   NOR2_X1 i_1_66 (.A1(n_1_857), .A2(n_267), .ZN(n_130));
   NOR2_X1 i_1_67 (.A1(n_1_858), .A2(n_267), .ZN(n_131));
   NOR3_X1 i_1_68 (.A1(counter[0]), .A2(n_267), .A3(n_1_657), .ZN(n_132));
   NOR2_X1 i_1_69 (.A1(n_1_794), .A2(n_1_6), .ZN(n_133));
   NOR2_X1 i_1_70 (.A1(n_1_793), .A2(n_1_6), .ZN(n_134));
   NOR2_X1 i_1_71 (.A1(n_1_792), .A2(n_1_6), .ZN(n_135));
   NOR2_X1 i_1_72 (.A1(n_1_791), .A2(n_1_6), .ZN(n_136));
   OAI21_X1 i_1_73 (.A(n_1_617), .B1(n_1_922), .B2(n_1_7), .ZN(n_1_6));
   AOI211_X1 i_1_74 (.A(reset), .B(resetReg), .C1(n_1_788), .C2(n_1_786), 
      .ZN(n_1_7));
   OAI21_X1 i_1_75 (.A(n_1_8), .B1(n_1_795), .B2(n_1_784), .ZN(n_137));
   NAND3_X1 i_1_76 (.A1(b[0]), .A2(a[0]), .A3(n_1_784), .ZN(n_1_8));
   OAI22_X1 i_1_77 (.A1(n_1_796), .A2(n_1_784), .B1(n_1_785), .B2(n_1_9), 
      .ZN(n_138));
   INV_X1 i_1_78 (.A(n_1_10), .ZN(n_1_9));
   OAI222_X1 i_1_79 (.A1(n_1_860), .A2(n_1_73), .B1(n_1_859), .B2(n_1_72), 
      .C1(n_1_891), .C2(n_1_71), .ZN(n_1_10));
   OAI22_X1 i_1_80 (.A1(n_1_797), .A2(n_1_784), .B1(n_1_785), .B2(n_1_11), 
      .ZN(n_139));
   INV_X1 i_1_81 (.A(n_1_12), .ZN(n_1_11));
   OAI222_X1 i_1_82 (.A1(n_1_861), .A2(n_1_73), .B1(n_1_891), .B2(n_1_72), 
      .C1(n_1_892), .C2(n_1_71), .ZN(n_1_12));
   OAI22_X1 i_1_83 (.A1(n_1_798), .A2(n_1_784), .B1(n_1_785), .B2(n_1_13), 
      .ZN(n_140));
   INV_X1 i_1_84 (.A(n_1_14), .ZN(n_1_13));
   OAI222_X1 i_1_85 (.A1(n_1_862), .A2(n_1_73), .B1(n_1_892), .B2(n_1_72), 
      .C1(n_1_893), .C2(n_1_71), .ZN(n_1_14));
   OAI22_X1 i_1_86 (.A1(n_1_799), .A2(n_1_784), .B1(n_1_785), .B2(n_1_15), 
      .ZN(n_141));
   INV_X1 i_1_87 (.A(n_1_16), .ZN(n_1_15));
   OAI222_X1 i_1_88 (.A1(n_1_863), .A2(n_1_73), .B1(n_1_893), .B2(n_1_72), 
      .C1(n_1_894), .C2(n_1_71), .ZN(n_1_16));
   OAI22_X1 i_1_89 (.A1(n_1_800), .A2(n_1_784), .B1(n_1_785), .B2(n_1_17), 
      .ZN(n_142));
   INV_X1 i_1_90 (.A(n_1_18), .ZN(n_1_17));
   OAI222_X1 i_1_91 (.A1(n_1_864), .A2(n_1_73), .B1(n_1_894), .B2(n_1_72), 
      .C1(n_1_895), .C2(n_1_71), .ZN(n_1_18));
   OAI22_X1 i_1_92 (.A1(n_1_801), .A2(n_1_784), .B1(n_1_785), .B2(n_1_19), 
      .ZN(n_143));
   INV_X1 i_1_93 (.A(n_1_20), .ZN(n_1_19));
   OAI222_X1 i_1_94 (.A1(n_1_865), .A2(n_1_73), .B1(n_1_895), .B2(n_1_72), 
      .C1(n_1_896), .C2(n_1_71), .ZN(n_1_20));
   OAI22_X1 i_1_95 (.A1(n_1_802), .A2(n_1_784), .B1(n_1_785), .B2(n_1_21), 
      .ZN(n_144));
   INV_X1 i_1_96 (.A(n_1_22), .ZN(n_1_21));
   OAI222_X1 i_1_97 (.A1(n_1_866), .A2(n_1_73), .B1(n_1_896), .B2(n_1_72), 
      .C1(n_1_897), .C2(n_1_71), .ZN(n_1_22));
   OAI22_X1 i_1_98 (.A1(n_1_803), .A2(n_1_784), .B1(n_1_785), .B2(n_1_23), 
      .ZN(n_145));
   INV_X1 i_1_99 (.A(n_1_24), .ZN(n_1_23));
   OAI222_X1 i_1_100 (.A1(n_1_867), .A2(n_1_73), .B1(n_1_897), .B2(n_1_72), 
      .C1(n_1_898), .C2(n_1_71), .ZN(n_1_24));
   OAI22_X1 i_1_101 (.A1(n_1_804), .A2(n_1_784), .B1(n_1_785), .B2(n_1_25), 
      .ZN(n_146));
   INV_X1 i_1_102 (.A(n_1_26), .ZN(n_1_25));
   OAI222_X1 i_1_103 (.A1(n_1_868), .A2(n_1_73), .B1(n_1_898), .B2(n_1_72), 
      .C1(n_1_899), .C2(n_1_71), .ZN(n_1_26));
   OAI22_X1 i_1_104 (.A1(n_1_805), .A2(n_1_784), .B1(n_1_785), .B2(n_1_27), 
      .ZN(n_147));
   INV_X1 i_1_105 (.A(n_1_28), .ZN(n_1_27));
   OAI222_X1 i_1_106 (.A1(n_1_869), .A2(n_1_73), .B1(n_1_899), .B2(n_1_72), 
      .C1(n_1_900), .C2(n_1_71), .ZN(n_1_28));
   OAI22_X1 i_1_107 (.A1(n_1_806), .A2(n_1_784), .B1(n_1_785), .B2(n_1_29), 
      .ZN(n_148));
   INV_X1 i_1_108 (.A(n_1_30), .ZN(n_1_29));
   OAI222_X1 i_1_109 (.A1(n_1_870), .A2(n_1_73), .B1(n_1_900), .B2(n_1_72), 
      .C1(n_1_901), .C2(n_1_71), .ZN(n_1_30));
   OAI22_X1 i_1_110 (.A1(n_1_807), .A2(n_1_784), .B1(n_1_785), .B2(n_1_31), 
      .ZN(n_149));
   INV_X1 i_1_111 (.A(n_1_32), .ZN(n_1_31));
   OAI222_X1 i_1_112 (.A1(n_1_871), .A2(n_1_73), .B1(n_1_901), .B2(n_1_72), 
      .C1(n_1_902), .C2(n_1_71), .ZN(n_1_32));
   OAI22_X1 i_1_113 (.A1(n_1_808), .A2(n_1_784), .B1(n_1_785), .B2(n_1_33), 
      .ZN(n_150));
   INV_X1 i_1_114 (.A(n_1_34), .ZN(n_1_33));
   OAI222_X1 i_1_115 (.A1(n_1_872), .A2(n_1_73), .B1(n_1_902), .B2(n_1_72), 
      .C1(n_1_903), .C2(n_1_71), .ZN(n_1_34));
   OAI22_X1 i_1_116 (.A1(n_1_809), .A2(n_1_784), .B1(n_1_785), .B2(n_1_35), 
      .ZN(n_151));
   INV_X1 i_1_117 (.A(n_1_36), .ZN(n_1_35));
   OAI222_X1 i_1_118 (.A1(n_1_873), .A2(n_1_73), .B1(n_1_903), .B2(n_1_72), 
      .C1(n_1_904), .C2(n_1_71), .ZN(n_1_36));
   OAI22_X1 i_1_119 (.A1(n_1_810), .A2(n_1_784), .B1(n_1_785), .B2(n_1_37), 
      .ZN(n_152));
   INV_X1 i_1_120 (.A(n_1_38), .ZN(n_1_37));
   OAI222_X1 i_1_121 (.A1(n_1_874), .A2(n_1_73), .B1(n_1_904), .B2(n_1_72), 
      .C1(n_1_905), .C2(n_1_71), .ZN(n_1_38));
   OAI22_X1 i_1_122 (.A1(n_1_811), .A2(n_1_784), .B1(n_1_785), .B2(n_1_39), 
      .ZN(n_153));
   INV_X1 i_1_123 (.A(n_1_40), .ZN(n_1_39));
   OAI222_X1 i_1_124 (.A1(n_1_875), .A2(n_1_73), .B1(n_1_905), .B2(n_1_72), 
      .C1(n_1_906), .C2(n_1_71), .ZN(n_1_40));
   OAI22_X1 i_1_125 (.A1(n_1_812), .A2(n_1_784), .B1(n_1_785), .B2(n_1_41), 
      .ZN(n_154));
   INV_X1 i_1_126 (.A(n_1_42), .ZN(n_1_41));
   OAI222_X1 i_1_127 (.A1(n_1_876), .A2(n_1_73), .B1(n_1_906), .B2(n_1_72), 
      .C1(n_1_907), .C2(n_1_71), .ZN(n_1_42));
   OAI22_X1 i_1_128 (.A1(n_1_813), .A2(n_1_784), .B1(n_1_785), .B2(n_1_43), 
      .ZN(n_155));
   INV_X1 i_1_129 (.A(n_1_44), .ZN(n_1_43));
   OAI222_X1 i_1_130 (.A1(n_1_877), .A2(n_1_73), .B1(n_1_907), .B2(n_1_72), 
      .C1(n_1_908), .C2(n_1_71), .ZN(n_1_44));
   OAI22_X1 i_1_131 (.A1(n_1_814), .A2(n_1_784), .B1(n_1_785), .B2(n_1_45), 
      .ZN(n_156));
   INV_X1 i_1_132 (.A(n_1_46), .ZN(n_1_45));
   OAI222_X1 i_1_133 (.A1(n_1_878), .A2(n_1_73), .B1(n_1_908), .B2(n_1_72), 
      .C1(n_1_909), .C2(n_1_71), .ZN(n_1_46));
   OAI22_X1 i_1_134 (.A1(n_1_815), .A2(n_1_784), .B1(n_1_785), .B2(n_1_47), 
      .ZN(n_157));
   INV_X1 i_1_135 (.A(n_1_48), .ZN(n_1_47));
   OAI222_X1 i_1_136 (.A1(n_1_879), .A2(n_1_73), .B1(n_1_909), .B2(n_1_72), 
      .C1(n_1_910), .C2(n_1_71), .ZN(n_1_48));
   OAI22_X1 i_1_137 (.A1(n_1_816), .A2(n_1_784), .B1(n_1_785), .B2(n_1_49), 
      .ZN(n_158));
   INV_X1 i_1_138 (.A(n_1_50), .ZN(n_1_49));
   OAI222_X1 i_1_139 (.A1(n_1_880), .A2(n_1_73), .B1(n_1_910), .B2(n_1_72), 
      .C1(n_1_911), .C2(n_1_71), .ZN(n_1_50));
   OAI22_X1 i_1_140 (.A1(n_1_817), .A2(n_1_784), .B1(n_1_785), .B2(n_1_51), 
      .ZN(n_159));
   INV_X1 i_1_141 (.A(n_1_52), .ZN(n_1_51));
   OAI222_X1 i_1_142 (.A1(n_1_881), .A2(n_1_73), .B1(n_1_911), .B2(n_1_72), 
      .C1(n_1_912), .C2(n_1_71), .ZN(n_1_52));
   OAI22_X1 i_1_143 (.A1(n_1_818), .A2(n_1_784), .B1(n_1_785), .B2(n_1_53), 
      .ZN(n_160));
   INV_X1 i_1_144 (.A(n_1_54), .ZN(n_1_53));
   OAI222_X1 i_1_145 (.A1(n_1_882), .A2(n_1_73), .B1(n_1_912), .B2(n_1_72), 
      .C1(n_1_913), .C2(n_1_71), .ZN(n_1_54));
   OAI22_X1 i_1_146 (.A1(n_1_819), .A2(n_1_784), .B1(n_1_785), .B2(n_1_55), 
      .ZN(n_161));
   INV_X1 i_1_147 (.A(n_1_56), .ZN(n_1_55));
   OAI222_X1 i_1_148 (.A1(n_1_883), .A2(n_1_73), .B1(n_1_913), .B2(n_1_72), 
      .C1(n_1_914), .C2(n_1_71), .ZN(n_1_56));
   OAI22_X1 i_1_149 (.A1(n_1_820), .A2(n_1_784), .B1(n_1_785), .B2(n_1_57), 
      .ZN(n_162));
   INV_X1 i_1_150 (.A(n_1_58), .ZN(n_1_57));
   OAI222_X1 i_1_151 (.A1(n_1_884), .A2(n_1_73), .B1(n_1_914), .B2(n_1_72), 
      .C1(n_1_915), .C2(n_1_71), .ZN(n_1_58));
   OAI22_X1 i_1_152 (.A1(n_1_821), .A2(n_1_784), .B1(n_1_785), .B2(n_1_59), 
      .ZN(n_163));
   INV_X1 i_1_153 (.A(n_1_60), .ZN(n_1_59));
   OAI222_X1 i_1_154 (.A1(n_1_885), .A2(n_1_73), .B1(n_1_915), .B2(n_1_72), 
      .C1(n_1_916), .C2(n_1_71), .ZN(n_1_60));
   OAI22_X1 i_1_155 (.A1(n_1_822), .A2(n_1_784), .B1(n_1_785), .B2(n_1_61), 
      .ZN(n_164));
   INV_X1 i_1_156 (.A(n_1_62), .ZN(n_1_61));
   OAI222_X1 i_1_157 (.A1(n_1_886), .A2(n_1_73), .B1(n_1_916), .B2(n_1_72), 
      .C1(n_1_917), .C2(n_1_71), .ZN(n_1_62));
   OAI22_X1 i_1_158 (.A1(n_1_823), .A2(n_1_784), .B1(n_1_785), .B2(n_1_63), 
      .ZN(n_165));
   INV_X1 i_1_159 (.A(n_1_64), .ZN(n_1_63));
   OAI222_X1 i_1_160 (.A1(n_1_887), .A2(n_1_73), .B1(n_1_917), .B2(n_1_72), 
      .C1(n_1_918), .C2(n_1_71), .ZN(n_1_64));
   OAI22_X1 i_1_161 (.A1(n_1_824), .A2(n_1_784), .B1(n_1_785), .B2(n_1_65), 
      .ZN(n_166));
   INV_X1 i_1_162 (.A(n_1_66), .ZN(n_1_65));
   OAI222_X1 i_1_163 (.A1(n_1_888), .A2(n_1_73), .B1(n_1_918), .B2(n_1_72), 
      .C1(n_1_919), .C2(n_1_71), .ZN(n_1_66));
   OAI22_X1 i_1_164 (.A1(n_1_825), .A2(n_1_784), .B1(n_1_785), .B2(n_1_67), 
      .ZN(n_167));
   INV_X1 i_1_165 (.A(n_1_68), .ZN(n_1_67));
   OAI222_X1 i_1_166 (.A1(n_1_889), .A2(n_1_73), .B1(n_1_919), .B2(n_1_72), 
      .C1(n_1_920), .C2(n_1_71), .ZN(n_1_68));
   OAI21_X1 i_1_167 (.A(n_1_69), .B1(n_1_826), .B2(n_1_784), .ZN(n_168));
   OAI21_X1 i_1_168 (.A(n_1_69), .B1(n_1_827), .B2(n_1_784), .ZN(n_169));
   OAI21_X1 i_1_169 (.A(n_1_69), .B1(n_1_828), .B2(n_1_784), .ZN(n_170));
   OAI21_X1 i_1_170 (.A(n_1_69), .B1(n_1_829), .B2(n_1_784), .ZN(n_171));
   OAI21_X1 i_1_171 (.A(n_1_69), .B1(n_1_830), .B2(n_1_784), .ZN(n_172));
   OAI21_X1 i_1_172 (.A(n_1_69), .B1(n_1_831), .B2(n_1_784), .ZN(n_173));
   OAI21_X1 i_1_173 (.A(n_1_69), .B1(n_1_832), .B2(n_1_784), .ZN(n_174));
   OAI21_X1 i_1_174 (.A(n_1_69), .B1(n_1_833), .B2(n_1_784), .ZN(n_175));
   OAI21_X1 i_1_175 (.A(n_1_69), .B1(n_1_834), .B2(n_1_784), .ZN(n_176));
   OAI21_X1 i_1_176 (.A(n_1_69), .B1(n_1_835), .B2(n_1_784), .ZN(n_177));
   OAI21_X1 i_1_177 (.A(n_1_69), .B1(n_1_836), .B2(n_1_784), .ZN(n_178));
   OAI21_X1 i_1_178 (.A(n_1_69), .B1(n_1_837), .B2(n_1_784), .ZN(n_179));
   OAI21_X1 i_1_179 (.A(n_1_69), .B1(n_1_838), .B2(n_1_784), .ZN(n_180));
   OAI21_X1 i_1_180 (.A(n_1_69), .B1(n_1_839), .B2(n_1_784), .ZN(n_181));
   OAI21_X1 i_1_181 (.A(n_1_69), .B1(n_1_840), .B2(n_1_784), .ZN(n_182));
   OAI21_X1 i_1_182 (.A(n_1_69), .B1(n_1_841), .B2(n_1_784), .ZN(n_183));
   OAI21_X1 i_1_183 (.A(n_1_69), .B1(n_1_842), .B2(n_1_784), .ZN(n_184));
   OAI21_X1 i_1_184 (.A(n_1_69), .B1(n_1_843), .B2(n_1_784), .ZN(n_185));
   OAI21_X1 i_1_185 (.A(n_1_69), .B1(n_1_844), .B2(n_1_784), .ZN(n_186));
   OAI21_X1 i_1_186 (.A(n_1_69), .B1(n_1_845), .B2(n_1_784), .ZN(n_187));
   OAI21_X1 i_1_187 (.A(n_1_69), .B1(n_1_846), .B2(n_1_784), .ZN(n_188));
   OAI21_X1 i_1_188 (.A(n_1_69), .B1(n_1_847), .B2(n_1_784), .ZN(n_189));
   OAI21_X1 i_1_189 (.A(n_1_69), .B1(n_1_848), .B2(n_1_784), .ZN(n_190));
   OAI21_X1 i_1_190 (.A(n_1_69), .B1(n_1_849), .B2(n_1_784), .ZN(n_191));
   OAI21_X1 i_1_191 (.A(n_1_69), .B1(n_1_850), .B2(n_1_784), .ZN(n_192));
   OAI21_X1 i_1_192 (.A(n_1_69), .B1(n_1_851), .B2(n_1_784), .ZN(n_193));
   OAI21_X1 i_1_193 (.A(n_1_69), .B1(n_1_852), .B2(n_1_784), .ZN(n_194));
   OAI21_X1 i_1_194 (.A(n_1_69), .B1(n_1_853), .B2(n_1_784), .ZN(n_195));
   OAI21_X1 i_1_195 (.A(n_1_69), .B1(n_1_854), .B2(n_1_784), .ZN(n_196));
   OAI21_X1 i_1_196 (.A(n_1_69), .B1(n_1_855), .B2(n_1_784), .ZN(n_197));
   OAI21_X1 i_1_197 (.A(n_1_69), .B1(n_1_856), .B2(n_1_784), .ZN(n_198));
   OAI21_X1 i_1_198 (.A(n_1_69), .B1(n_1_857), .B2(n_1_784), .ZN(n_199));
   OAI21_X1 i_1_199 (.A(n_1_69), .B1(n_1_858), .B2(n_1_784), .ZN(n_200));
   NAND2_X1 i_1_200 (.A1(n_1_784), .A2(n_1_70), .ZN(n_1_69));
   OAI222_X1 i_1_201 (.A1(n_1_920), .A2(n_1_72), .B1(n_1_921), .B2(n_1_71), 
      .C1(n_1_890), .C2(n_1_73), .ZN(n_1_70));
   NAND2_X1 i_1_202 (.A1(b[1]), .A2(b[0]), .ZN(n_1_71));
   NAND2_X1 i_1_203 (.A1(b[1]), .A2(n_1_923), .ZN(n_1_72));
   NAND2_X1 i_1_204 (.A1(n_1_924), .A2(b[0]), .ZN(n_1_73));
   NOR2_X1 i_1_205 (.A1(n_1_785), .A2(n_1_584), .ZN(n_201));
   NOR2_X1 i_1_206 (.A1(n_1_785), .A2(n_1_674), .ZN(n_202));
   OAI22_X1 i_1_207 (.A1(n_1_696), .A2(n_1_584), .B1(n_1_785), .B2(n_1_531), 
      .ZN(n_203));
   OAI22_X1 i_1_208 (.A1(n_1_696), .A2(n_1_674), .B1(n_1_785), .B2(n_1_678), 
      .ZN(n_204));
   OAI222_X1 i_1_209 (.A1(n_1_696), .A2(n_1_531), .B1(n_1_584), .B2(n_1_224), 
      .C1(n_1_785), .C2(n_1_575), .ZN(n_205));
   OAI222_X1 i_1_210 (.A1(n_1_674), .A2(n_1_224), .B1(n_1_696), .B2(n_1_678), 
      .C1(n_1_785), .C2(n_1_600), .ZN(n_206));
   OAI221_X1 i_1_211 (.A(n_1_74), .B1(n_1_785), .B2(n_1_578), .C1(n_1_584), 
      .C2(n_1_247), .ZN(n_207));
   AOI22_X1 i_1_212 (.A1(n_1_697), .A2(n_1_576), .B1(n_1_532), .B2(n_1_225), 
      .ZN(n_1_74));
   OAI221_X1 i_1_213 (.A(n_1_75), .B1(n_1_674), .B2(n_1_247), .C1(n_1_678), 
      .C2(n_1_224), .ZN(n_208));
   AOI22_X1 i_1_214 (.A1(n_1_784), .A2(n_1_665), .B1(n_1_697), .B2(n_1_601), 
      .ZN(n_1_75));
   OAI221_X1 i_1_215 (.A(n_1_76), .B1(n_1_575), .B2(n_1_224), .C1(n_1_692), 
      .C2(n_1_584), .ZN(n_209));
   AOI222_X1 i_1_216 (.A1(n_1_784), .A2(n_1_535), .B1(n_1_697), .B2(n_1_579), 
      .C1(n_1_532), .C2(n_1_248), .ZN(n_1_76));
   OAI221_X1 i_1_217 (.A(n_1_77), .B1(n_1_600), .B2(n_1_224), .C1(n_1_785), 
      .C2(n_1_649), .ZN(n_210));
   AOI21_X1 i_1_218 (.A(n_1_78), .B1(n_1_697), .B2(n_1_665), .ZN(n_1_77));
   OAI22_X1 i_1_219 (.A1(n_1_692), .A2(n_1_674), .B1(n_1_678), .B2(n_1_247), 
      .ZN(n_1_78));
   OAI221_X1 i_1_220 (.A(n_1_79), .B1(n_1_785), .B2(n_1_547), .C1(n_1_707), 
      .C2(n_1_584), .ZN(n_211));
   AOI221_X1 i_1_221 (.A(n_1_80), .B1(n_1_576), .B2(n_1_248), .C1(n_1_697), 
      .C2(n_1_535), .ZN(n_1_79));
   OAI22_X1 i_1_222 (.A1(n_1_692), .A2(n_1_531), .B1(n_1_578), .B2(n_1_224), 
      .ZN(n_1_80));
   OAI221_X1 i_1_223 (.A(n_1_81), .B1(n_1_707), .B2(n_1_674), .C1(n_1_600), 
      .C2(n_1_247), .ZN(n_212));
   AOI221_X1 i_1_224 (.A(n_1_82), .B1(n_1_665), .B2(n_1_225), .C1(n_1_697), 
      .C2(n_1_650), .ZN(n_1_81));
   OAI22_X1 i_1_225 (.A1(n_1_692), .A2(n_1_678), .B1(n_1_785), .B2(n_1_625), 
      .ZN(n_1_82));
   OAI211_X1 i_1_226 (.A(n_1_85), .B(n_1_83), .C1(n_1_534), .C2(n_1_224), 
      .ZN(n_213));
   AOI221_X1 i_1_227 (.A(n_1_84), .B1(n_1_697), .B2(n_1_548), .C1(n_1_579), 
      .C2(n_1_248), .ZN(n_1_83));
   OAI22_X1 i_1_228 (.A1(n_1_785), .A2(n_1_541), .B1(n_1_713), .B2(n_1_584), 
      .ZN(n_1_84));
   INV_X1 i_1_229 (.A(n_1_86), .ZN(n_1_85));
   OAI22_X1 i_1_230 (.A1(n_1_692), .A2(n_1_575), .B1(n_1_707), .B2(n_1_531), 
      .ZN(n_1_86));
   OAI211_X1 i_1_231 (.A(n_1_89), .B(n_1_87), .C1(n_1_696), .C2(n_1_625), 
      .ZN(n_214));
   AOI221_X1 i_1_232 (.A(n_1_88), .B1(n_1_650), .B2(n_1_225), .C1(n_1_708), 
      .C2(n_1_679), .ZN(n_1_87));
   OAI22_X1 i_1_233 (.A1(n_1_692), .A2(n_1_600), .B1(n_1_664), .B2(n_1_247), 
      .ZN(n_1_88));
   AOI22_X1 i_1_234 (.A1(n_1_712), .A2(n_1_675), .B1(n_1_784), .B2(n_1_685), 
      .ZN(n_1_89));
   OR3_X1 i_1_235 (.A1(n_1_93), .A2(n_1_92), .A3(n_1_90), .ZN(n_215));
   OAI221_X1 i_1_236 (.A(n_1_91), .B1(n_1_713), .B2(n_1_531), .C1(n_1_584), 
      .C2(n_1_486), .ZN(n_1_90));
   AOI22_X1 i_1_237 (.A1(n_1_784), .A2(n_1_582), .B1(n_1_708), .B2(n_1_576), 
      .ZN(n_1_91));
   OAI22_X1 i_1_238 (.A1(n_1_534), .A2(n_1_247), .B1(n_1_692), .B2(n_1_578), 
      .ZN(n_1_92));
   OAI22_X1 i_1_239 (.A1(n_1_547), .A2(n_1_224), .B1(n_1_696), .B2(n_1_541), 
      .ZN(n_1_93));
   OR3_X1 i_1_240 (.A1(n_1_97), .A2(n_1_96), .A3(n_1_94), .ZN(n_216));
   OAI221_X1 i_1_241 (.A(n_1_95), .B1(n_1_692), .B2(n_1_664), .C1(n_1_707), 
      .C2(n_1_600), .ZN(n_1_94));
   AOI22_X1 i_1_242 (.A1(n_1_675), .A2(n_1_487), .B1(n_1_712), .B2(n_1_679), 
      .ZN(n_1_95));
   OAI22_X1 i_1_243 (.A1(n_1_785), .A2(n_1_629), .B1(n_1_696), .B2(n_1_684), 
      .ZN(n_1_96));
   OAI22_X1 i_1_244 (.A1(n_1_649), .A2(n_1_247), .B1(n_1_625), .B2(n_1_224), 
      .ZN(n_1_97));
   INV_X1 i_1_245 (.A(n_1_98), .ZN(n_217));
   AOI211_X1 i_1_246 (.A(n_1_102), .B(n_1_99), .C1(n_1_542), .C2(n_1_225), 
      .ZN(n_1_98));
   OAI221_X1 i_1_247 (.A(n_1_100), .B1(n_1_531), .B2(n_1_486), .C1(n_1_704), 
      .C2(n_1_584), .ZN(n_1_99));
   AOI221_X1 i_1_248 (.A(n_1_101), .B1(n_1_712), .B2(n_1_576), .C1(n_1_784), 
      .C2(n_1_551), .ZN(n_1_100));
   OAI22_X1 i_1_249 (.A1(n_1_696), .A2(n_1_581), .B1(n_1_547), .B2(n_1_247), 
      .ZN(n_1_101));
   OAI22_X1 i_1_250 (.A1(n_1_692), .A2(n_1_534), .B1(n_1_707), .B2(n_1_578), 
      .ZN(n_1_102));
   INV_X1 i_1_251 (.A(n_1_103), .ZN(n_218));
   AOI211_X1 i_1_252 (.A(n_1_107), .B(n_1_104), .C1(n_1_708), .C2(n_1_665), 
      .ZN(n_1_103));
   OAI221_X1 i_1_253 (.A(n_1_105), .B1(n_1_684), .B2(n_1_224), .C1(n_1_713), 
      .C2(n_1_600), .ZN(n_1_104));
   AOI221_X1 i_1_254 (.A(n_1_106), .B1(n_1_626), .B2(n_1_248), .C1(n_1_679), 
      .C2(n_1_487), .ZN(n_1_105));
   OAI22_X1 i_1_255 (.A1(n_1_704), .A2(n_1_674), .B1(n_1_696), .B2(n_1_629), 
      .ZN(n_1_106));
   OAI22_X1 i_1_256 (.A1(n_1_785), .A2(n_1_670), .B1(n_1_692), .B2(n_1_649), 
      .ZN(n_1_107));
   OR3_X1 i_1_257 (.A1(n_1_112), .A2(n_1_111), .A3(n_1_108), .ZN(n_219));
   OAI221_X1 i_1_258 (.A(n_1_109), .B1(n_1_701), .B2(n_1_584), .C1(n_1_696), 
      .C2(n_1_550), .ZN(n_1_108));
   AOI221_X1 i_1_259 (.A(n_1_110), .B1(n_1_708), .B2(n_1_535), .C1(n_1_542), 
      .C2(n_1_248), .ZN(n_1_109));
   OAI22_X1 i_1_260 (.A1(n_1_581), .A2(n_1_224), .B1(n_1_692), .B2(n_1_547), 
      .ZN(n_1_110));
   OAI22_X1 i_1_261 (.A1(n_1_713), .A2(n_1_578), .B1(n_1_785), .B2(n_1_566), 
      .ZN(n_1_111));
   OAI22_X1 i_1_262 (.A1(n_1_575), .A2(n_1_486), .B1(n_1_704), .B2(n_1_531), 
      .ZN(n_1_112));
   OR3_X1 i_1_263 (.A1(n_1_117), .A2(n_1_116), .A3(n_1_113), .ZN(n_220));
   OAI221_X1 i_1_264 (.A(n_1_114), .B1(n_1_785), .B2(n_1_596), .C1(n_1_696), 
      .C2(n_1_670), .ZN(n_1_113));
   AOI221_X1 i_1_265 (.A(n_1_115), .B1(n_1_712), .B2(n_1_665), .C1(n_1_708), 
      .C2(n_1_650), .ZN(n_1_114));
   OAI22_X1 i_1_266 (.A1(n_1_692), .A2(n_1_625), .B1(n_1_701), .B2(n_1_674), 
      .ZN(n_1_115));
   OAI22_X1 i_1_267 (.A1(n_1_629), .A2(n_1_224), .B1(n_1_704), .B2(n_1_678), 
      .ZN(n_1_116));
   OAI22_X1 i_1_268 (.A1(n_1_684), .A2(n_1_247), .B1(n_1_600), .B2(n_1_486), 
      .ZN(n_1_117));
   OR4_X1 i_1_269 (.A1(n_1_119), .A2(n_1_118), .A3(n_1_120), .A4(n_1_122), 
      .ZN(n_221));
   OAI22_X1 i_1_270 (.A1(n_1_550), .A2(n_1_224), .B1(n_1_581), .B2(n_1_247), 
      .ZN(n_1_118));
   OAI22_X1 i_1_271 (.A1(n_1_696), .A2(n_1_566), .B1(n_1_724), .B2(n_1_584), 
      .ZN(n_1_119));
   OAI221_X1 i_1_272 (.A(n_1_121), .B1(n_1_713), .B2(n_1_534), .C1(n_1_785), 
      .C2(n_1_538), .ZN(n_1_120));
   AOI22_X1 i_1_273 (.A1(n_1_708), .A2(n_1_548), .B1(n_1_579), .B2(n_1_487), 
      .ZN(n_1_121));
   OAI222_X1 i_1_274 (.A1(n_1_704), .A2(n_1_575), .B1(n_1_692), .B2(n_1_541), 
      .C1(n_1_701), .C2(n_1_531), .ZN(n_1_122));
   OR4_X1 i_1_275 (.A1(n_1_124), .A2(n_1_123), .A3(n_1_125), .A4(n_1_128), 
      .ZN(n_222));
   OAI22_X1 i_1_276 (.A1(n_1_724), .A2(n_1_674), .B1(n_1_713), .B2(n_1_649), 
      .ZN(n_1_123));
   OAI22_X1 i_1_277 (.A1(n_1_785), .A2(n_1_609), .B1(n_1_664), .B2(n_1_486), 
      .ZN(n_1_124));
   OAI221_X1 i_1_278 (.A(n_1_126), .B1(n_1_701), .B2(n_1_678), .C1(n_1_707), 
      .C2(n_1_625), .ZN(n_1_125));
   INV_X1 i_1_279 (.A(n_1_127), .ZN(n_1_126));
   OAI22_X1 i_1_280 (.A1(n_1_629), .A2(n_1_247), .B1(n_1_692), .B2(n_1_684), 
      .ZN(n_1_127));
   OAI222_X1 i_1_281 (.A1(n_1_704), .A2(n_1_600), .B1(n_1_670), .B2(n_1_224), 
      .C1(n_1_696), .C2(n_1_596), .ZN(n_1_128));
   OR4_X1 i_1_282 (.A1(n_1_130), .A2(n_1_129), .A3(n_1_131), .A4(n_1_134), 
      .ZN(n_223));
   OAI22_X1 i_1_283 (.A1(n_1_550), .A2(n_1_247), .B1(n_1_713), .B2(n_1_547), 
      .ZN(n_1_129));
   OAI22_X1 i_1_284 (.A1(n_1_724), .A2(n_1_531), .B1(n_1_661), .B2(n_1_584), 
      .ZN(n_1_130));
   OAI221_X1 i_1_285 (.A(n_1_132), .B1(n_1_704), .B2(n_1_578), .C1(n_1_785), 
      .C2(n_1_553), .ZN(n_1_131));
   INV_X1 i_1_286 (.A(n_1_133), .ZN(n_1_132));
   OAI22_X1 i_1_287 (.A1(n_1_707), .A2(n_1_541), .B1(n_1_692), .B2(n_1_581), 
      .ZN(n_1_133));
   OAI221_X1 i_1_288 (.A(n_1_135), .B1(n_1_534), .B2(n_1_486), .C1(n_1_701), 
      .C2(n_1_575), .ZN(n_1_134));
   AOI22_X1 i_1_289 (.A1(n_1_567), .A2(n_1_225), .B1(n_1_697), .B2(n_1_539), 
      .ZN(n_1_135));
   OR4_X1 i_1_290 (.A1(n_1_137), .A2(n_1_136), .A3(n_1_138), .A4(n_1_141), 
      .ZN(n_224));
   OAI22_X1 i_1_291 (.A1(n_1_596), .A2(n_1_224), .B1(n_1_707), .B2(n_1_684), 
      .ZN(n_1_136));
   OAI22_X1 i_1_292 (.A1(n_1_692), .A2(n_1_629), .B1(n_1_674), .B2(n_1_661), 
      .ZN(n_1_137));
   OAI221_X1 i_1_293 (.A(n_1_139), .B1(n_1_670), .B2(n_1_247), .C1(n_1_785), 
      .C2(n_1_605), .ZN(n_1_138));
   INV_X1 i_1_294 (.A(n_1_140), .ZN(n_1_139));
   OAI22_X1 i_1_295 (.A1(n_1_701), .A2(n_1_600), .B1(n_1_704), .B2(n_1_664), 
      .ZN(n_1_140));
   OAI221_X1 i_1_296 (.A(n_1_142), .B1(n_1_649), .B2(n_1_486), .C1(n_1_713), 
      .C2(n_1_625), .ZN(n_1_141));
   AOI22_X1 i_1_297 (.A1(n_1_697), .A2(n_1_610), .B1(n_1_725), .B2(n_1_679), 
      .ZN(n_1_142));
   OR3_X1 i_1_298 (.A1(n_1_145), .A2(n_1_143), .A3(n_1_146), .ZN(n_225));
   OAI221_X1 i_1_299 (.A(n_1_144), .B1(n_1_692), .B2(n_1_550), .C1(n_1_538), 
      .C2(n_1_224), .ZN(n_1_143));
   AOI22_X1 i_1_300 (.A1(n_1_708), .A2(n_1_582), .B1(n_1_784), .B2(n_1_557), 
      .ZN(n_1_144));
   OAI222_X1 i_1_301 (.A1(n_1_701), .A2(n_1_578), .B1(n_1_724), .B2(n_1_575), 
      .C1(n_1_713), .C2(n_1_541), .ZN(n_1_145));
   OAI221_X1 i_1_302 (.A(n_1_147), .B1(n_1_704), .B2(n_1_534), .C1(n_1_645), 
      .C2(n_1_584), .ZN(n_1_146));
   AOI221_X1 i_1_303 (.A(n_1_148), .B1(n_1_567), .B2(n_1_248), .C1(n_1_662), 
      .C2(n_1_532), .ZN(n_1_147));
   OAI22_X1 i_1_304 (.A1(n_1_547), .A2(n_1_486), .B1(n_1_696), .B2(n_1_553), 
      .ZN(n_1_148));
   OR4_X1 i_1_305 (.A1(n_1_150), .A2(n_1_149), .A3(n_1_151), .A4(n_1_152), 
      .ZN(n_226));
   OAI22_X1 i_1_306 (.A1(n_1_713), .A2(n_1_684), .B1(n_1_609), .B2(n_1_224), 
      .ZN(n_1_149));
   OAI22_X1 i_1_307 (.A1(n_1_596), .A2(n_1_247), .B1(n_1_707), .B2(n_1_629), 
      .ZN(n_1_150));
   OAI222_X1 i_1_308 (.A1(n_1_704), .A2(n_1_649), .B1(n_1_701), .B2(n_1_664), 
      .C1(n_1_678), .C2(n_1_661), .ZN(n_1_151));
   OAI221_X1 i_1_309 (.A(n_1_153), .B1(n_1_785), .B2(n_1_637), .C1(n_1_696), 
      .C2(n_1_605), .ZN(n_1_152));
   AOI221_X1 i_1_310 (.A(n_1_154), .B1(n_1_626), .B2(n_1_487), .C1(n_1_725), 
      .C2(n_1_601), .ZN(n_1_153));
   OAI22_X1 i_1_311 (.A1(n_1_674), .A2(n_1_645), .B1(n_1_692), .B2(n_1_670), 
      .ZN(n_1_154));
   OR4_X1 i_1_312 (.A1(n_1_156), .A2(n_1_155), .A3(n_1_157), .A4(n_1_159), 
      .ZN(n_227));
   OAI22_X1 i_1_313 (.A1(n_1_538), .A2(n_1_247), .B1(n_1_645), .B2(n_1_531), 
      .ZN(n_1_155));
   OAI22_X1 i_1_314 (.A1(n_1_724), .A2(n_1_578), .B1(n_1_704), .B2(n_1_547), 
      .ZN(n_1_156));
   OAI221_X1 i_1_315 (.A(n_1_158), .B1(n_1_692), .B2(n_1_566), .C1(n_1_785), 
      .C2(n_1_560), .ZN(n_1_157));
   AOI22_X1 i_1_316 (.A1(n_1_542), .A2(n_1_487), .B1(n_1_662), .B2(n_1_576), 
      .ZN(n_1_158));
   OAI221_X1 i_1_317 (.A(n_1_160), .B1(n_1_701), .B2(n_1_534), .C1(n_1_647), 
      .C2(n_1_584), .ZN(n_1_159));
   AOI221_X1 i_1_318 (.A(n_1_161), .B1(n_1_554), .B2(n_1_225), .C1(n_1_712), 
      .C2(n_1_582), .ZN(n_1_160));
   OAI22_X1 i_1_319 (.A1(n_1_696), .A2(n_1_556), .B1(n_1_707), .B2(n_1_550), 
      .ZN(n_1_161));
   OR4_X1 i_1_320 (.A1(n_1_163), .A2(n_1_162), .A3(n_1_164), .A4(n_1_166), 
      .ZN(n_228));
   OAI22_X1 i_1_321 (.A1(n_1_605), .A2(n_1_224), .B1(n_1_678), .B2(n_1_645), 
      .ZN(n_1_162));
   OAI22_X1 i_1_322 (.A1(n_1_684), .A2(n_1_486), .B1(n_1_609), .B2(n_1_247), 
      .ZN(n_1_163));
   OAI221_X1 i_1_323 (.A(n_1_165), .B1(n_1_692), .B2(n_1_596), .C1(n_1_707), 
      .C2(n_1_670), .ZN(n_1_164));
   AOI22_X1 i_1_324 (.A1(n_1_662), .A2(n_1_601), .B1(n_1_675), .B2(n_1_648), 
      .ZN(n_1_165));
   OAI221_X1 i_1_325 (.A(n_1_167), .B1(n_1_704), .B2(n_1_625), .C1(n_1_701), 
      .C2(n_1_649), .ZN(n_1_166));
   AOI221_X1 i_1_326 (.A(n_1_168), .B1(n_1_784), .B2(n_1_619), .C1(n_1_697), 
      .C2(n_1_638), .ZN(n_1_167));
   OAI22_X1 i_1_327 (.A1(n_1_724), .A2(n_1_664), .B1(n_1_713), .B2(n_1_629), 
      .ZN(n_1_168));
   OR4_X1 i_1_328 (.A1(n_1_174), .A2(n_1_172), .A3(n_1_171), .A4(n_1_169), 
      .ZN(n_229));
   OAI221_X1 i_1_329 (.A(n_1_170), .B1(n_1_645), .B2(n_1_575), .C1(n_1_696), 
      .C2(n_1_560), .ZN(n_1_169));
   AOI22_X1 i_1_330 (.A1(n_1_784), .A2(n_1_573), .B1(n_1_648), .B2(n_1_532), 
      .ZN(n_1_170));
   OAI222_X1 i_1_331 (.A1(n_1_556), .A2(n_1_224), .B1(n_1_553), .B2(n_1_247), 
      .C1(n_1_704), .C2(n_1_541), .ZN(n_1_171));
   OAI221_X1 i_1_332 (.A(n_1_173), .B1(n_1_713), .B2(n_1_550), .C1(n_1_584), 
      .C2(n_1_516), .ZN(n_1_172));
   AOI22_X1 i_1_333 (.A1(n_1_708), .A2(n_1_567), .B1(n_1_582), .B2(n_1_487), 
      .ZN(n_1_173));
   OAI221_X1 i_1_334 (.A(n_1_175), .B1(n_1_701), .B2(n_1_547), .C1(n_1_661), 
      .C2(n_1_578), .ZN(n_1_174));
   INV_X1 i_1_335 (.A(n_1_176), .ZN(n_1_175));
   OAI22_X1 i_1_336 (.A1(n_1_724), .A2(n_1_534), .B1(n_1_692), .B2(n_1_538), 
      .ZN(n_1_176));
   OR4_X1 i_1_337 (.A1(n_1_182), .A2(n_1_180), .A3(n_1_179), .A4(n_1_177), 
      .ZN(n_230));
   OAI221_X1 i_1_338 (.A(n_1_178), .B1(n_1_696), .B2(n_1_618), .C1(n_1_724), 
      .C2(n_1_649), .ZN(n_1_177));
   AOI22_X1 i_1_339 (.A1(n_1_679), .A2(n_1_648), .B1(n_1_630), .B2(n_1_487), 
      .ZN(n_1_178));
   OAI222_X1 i_1_340 (.A1(n_1_713), .A2(n_1_670), .B1(n_1_704), .B2(n_1_684), 
      .C1(n_1_785), .C2(n_1_653), .ZN(n_1_179));
   OAI221_X1 i_1_341 (.A(n_1_181), .B1(n_1_707), .B2(n_1_596), .C1(n_1_701), 
      .C2(n_1_625), .ZN(n_1_180));
   AOI22_X1 i_1_342 (.A1(n_1_606), .A2(n_1_248), .B1(n_1_638), .B2(n_1_225), 
      .ZN(n_1_181));
   OAI221_X1 i_1_343 (.A(n_1_183), .B1(n_1_645), .B2(n_1_600), .C1(n_1_692), 
      .C2(n_1_609), .ZN(n_1_182));
   AOI22_X1 i_1_344 (.A1(n_1_675), .A2(n_1_517), .B1(n_1_665), .B2(n_1_662), 
      .ZN(n_1_183));
   OR4_X1 i_1_345 (.A1(n_1_191), .A2(n_1_189), .A3(n_1_186), .A4(n_1_184), 
      .ZN(n_231));
   OAI221_X1 i_1_346 (.A(n_1_185), .B1(n_1_696), .B2(n_1_572), .C1(n_1_661), 
      .C2(n_1_534), .ZN(n_1_184));
   AOI22_X1 i_1_347 (.A1(n_1_557), .A2(n_1_248), .B1(n_1_725), .B2(n_1_548), 
      .ZN(n_1_185));
   OAI221_X1 i_1_348 (.A(n_1_187), .B1(n_1_550), .B2(n_1_486), .C1(n_1_785), 
      .C2(n_1_563), .ZN(n_1_186));
   INV_X1 i_1_349 (.A(n_1_188), .ZN(n_1_187));
   OAI22_X1 i_1_350 (.A1(n_1_692), .A2(n_1_553), .B1(n_1_704), .B2(n_1_581), 
      .ZN(n_1_188));
   OAI221_X1 i_1_351 (.A(n_1_190), .B1(n_1_645), .B2(n_1_578), .C1(n_1_584), 
      .C2(n_1_504), .ZN(n_1_189));
   AOI22_X1 i_1_352 (.A1(n_1_561), .A2(n_1_225), .B1(n_1_712), .B2(n_1_567), 
      .ZN(n_1_190));
   OAI221_X1 i_1_353 (.A(n_1_192), .B1(n_1_531), .B2(n_1_516), .C1(n_1_701), 
      .C2(n_1_541), .ZN(n_1_191));
   AOI22_X1 i_1_354 (.A1(n_1_708), .A2(n_1_539), .B1(n_1_648), .B2(n_1_576), 
      .ZN(n_1_192));
   OR4_X1 i_1_355 (.A1(n_1_199), .A2(n_1_197), .A3(n_1_195), .A4(n_1_193), 
      .ZN(n_232));
   OAI221_X1 i_1_356 (.A(n_1_194), .B1(n_1_647), .B2(n_1_600), .C1(n_1_724), 
      .C2(n_1_625), .ZN(n_1_193));
   AOI22_X1 i_1_357 (.A1(n_1_665), .A2(n_1_646), .B1(n_1_638), .B2(n_1_248), 
      .ZN(n_1_194));
   OAI221_X1 i_1_358 (.A(n_1_196), .B1(n_1_692), .B2(n_1_605), .C1(n_1_704), 
      .C2(n_1_629), .ZN(n_1_195));
   AOI22_X1 i_1_359 (.A1(n_1_712), .A2(n_1_597), .B1(n_1_708), .B2(n_1_610), 
      .ZN(n_1_196));
   OAI221_X1 i_1_360 (.A(n_1_198), .B1(n_1_618), .B2(n_1_224), .C1(n_1_696), 
      .C2(n_1_653), .ZN(n_1_197));
   AOI21_X1 i_1_361 (.A(n_1_699), .B1(n_1_662), .B2(n_1_650), .ZN(n_1_198));
   OAI221_X1 i_1_362 (.A(n_1_200), .B1(n_1_678), .B2(n_1_516), .C1(n_1_674), 
      .C2(n_1_504), .ZN(n_1_199));
   AOI22_X1 i_1_363 (.A1(n_1_671), .A2(n_1_487), .B1(n_1_702), .B2(n_1_685), 
      .ZN(n_1_200));
   OR4_X1 i_1_364 (.A1(n_1_203), .A2(n_1_201), .A3(n_1_205), .A4(n_1_206), 
      .ZN(n_233));
   OAI221_X1 i_1_365 (.A(n_1_202), .B1(n_1_566), .B2(n_1_486), .C1(n_1_531), 
      .C2(n_1_504), .ZN(n_1_201));
   AOI22_X1 i_1_366 (.A1(n_1_725), .A2(n_1_542), .B1(n_1_662), .B2(n_1_548), 
      .ZN(n_1_202));
   OAI221_X1 i_1_367 (.A(n_1_204), .B1(n_1_575), .B2(n_1_516), .C1(n_1_713), 
      .C2(n_1_538), .ZN(n_1_203));
   AOI22_X1 i_1_368 (.A1(n_1_648), .A2(n_1_579), .B1(n_1_573), .B2(n_1_225), 
      .ZN(n_1_204));
   OAI222_X1 i_1_369 (.A1(n_1_707), .A2(n_1_553), .B1(n_1_645), .B2(n_1_534), 
      .C1(n_1_704), .C2(n_1_550), .ZN(n_1_205));
   OAI211_X1 i_1_370 (.A(n_1_698), .B(n_1_207), .C1(n_1_617), .C2(n_1_584), 
      .ZN(n_1_206));
   AOI221_X1 i_1_371 (.A(n_1_208), .B1(n_1_561), .B2(n_1_248), .C1(n_1_702), 
      .C2(n_1_582), .ZN(n_1_207));
   OAI22_X1 i_1_372 (.A1(n_1_696), .A2(n_1_563), .B1(n_1_692), .B2(n_1_556), 
      .ZN(n_1_208));
   OR3_X1 i_1_373 (.A1(n_1_693), .A2(n_1_215), .A3(n_1_209), .ZN(n_234));
   OR4_X1 i_1_374 (.A1(n_1_211), .A2(n_1_210), .A3(n_1_212), .A4(n_1_214), 
      .ZN(n_1_209));
   OAI22_X1 i_1_375 (.A1(n_1_692), .A2(n_1_637), .B1(n_1_704), .B2(n_1_670), 
      .ZN(n_1_210));
   OAI22_X1 i_1_376 (.A1(n_1_596), .A2(n_1_486), .B1(n_1_713), .B2(n_1_609), 
      .ZN(n_1_211));
   OAI221_X1 i_1_377 (.A(n_1_213), .B1(n_1_678), .B2(n_1_504), .C1(n_1_618), 
      .C2(n_1_247), .ZN(n_1_212));
   AOI22_X1 i_1_378 (.A1(n_1_654), .A2(n_1_225), .B1(n_1_725), .B2(n_1_685), 
      .ZN(n_1_213));
   OAI222_X1 i_1_379 (.A1(n_1_707), .A2(n_1_605), .B1(n_1_674), .B2(n_1_617), 
      .C1(n_1_649), .C2(n_1_645), .ZN(n_1_214));
   OAI221_X1 i_1_380 (.A(n_1_216), .B1(n_1_701), .B2(n_1_629), .C1(n_1_600), 
      .C2(n_1_516), .ZN(n_1_215));
   AOI22_X1 i_1_381 (.A1(n_1_665), .A2(n_1_648), .B1(n_1_662), .B2(n_1_626), 
      .ZN(n_1_216));
   OR4_X1 i_1_382 (.A1(n_1_227), .A2(n_1_226), .A3(n_1_693), .A4(n_1_217), 
      .ZN(n_235));
   OR4_X1 i_1_383 (.A1(n_1_221), .A2(n_1_220), .A3(n_1_218), .A4(n_1_222), 
      .ZN(n_1_217));
   OAI221_X1 i_1_384 (.A(n_1_219), .B1(n_1_578), .B2(n_1_516), .C1(n_1_575), 
      .C2(n_1_504), .ZN(n_1_218));
   AOI22_X1 i_1_385 (.A1(n_1_616), .A2(n_1_532), .B1(n_1_662), .B2(n_1_542), 
      .ZN(n_1_219));
   OAI22_X1 i_1_386 (.A1(n_1_704), .A2(n_1_566), .B1(n_1_692), .B2(n_1_560), 
      .ZN(n_1_220));
   OAI22_X1 i_1_387 (.A1(n_1_538), .A2(n_1_486), .B1(n_1_645), .B2(n_1_547), 
      .ZN(n_1_221));
   OAI221_X1 i_1_388 (.A(n_1_223), .B1(n_1_707), .B2(n_1_556), .C1(n_1_724), 
      .C2(n_1_581), .ZN(n_1_222));
   AOI22_X1 i_1_389 (.A1(n_1_564), .A2(n_1_225), .B1(n_1_702), .B2(n_1_551), 
      .ZN(n_1_223));
   INV_X1 i_1_390 (.A(n_1_225), .ZN(n_1_224));
   NOR2_X1 i_1_391 (.A1(n_1_727), .A2(n_1_722), .ZN(n_1_225));
   OAI22_X1 i_1_392 (.A1(n_1_713), .A2(n_1_553), .B1(n_1_647), .B2(n_1_534), 
      .ZN(n_1_226));
   OAI22_X1 i_1_393 (.A1(n_1_572), .A2(n_1_247), .B1(n_1_656), .B2(n_1_584), 
      .ZN(n_1_227));
   OR4_X1 i_1_394 (.A1(n_1_234), .A2(n_1_232), .A3(n_1_242), .A4(n_1_228), 
      .ZN(n_236));
   OAI211_X1 i_1_395 (.A(n_1_231), .B(n_1_229), .C1(n_1_707), .C2(n_1_637), 
      .ZN(n_1_228));
   AOI221_X1 i_1_396 (.A(n_1_230), .B1(n_1_610), .B2(n_1_487), .C1(n_1_601), 
      .C2(n_1_505), .ZN(n_1_229));
   OAI22_X1 i_1_397 (.A1(n_1_649), .A2(n_1_647), .B1(n_1_692), .B2(n_1_618), 
      .ZN(n_1_230));
   AOI22_X1 i_1_398 (.A1(n_1_646), .A2(n_1_626), .B1(n_1_685), .B2(n_1_662), 
      .ZN(n_1_231));
   OAI221_X1 i_1_399 (.A(n_1_233), .B1(n_1_674), .B2(n_1_656), .C1(n_1_701), 
      .C2(n_1_670), .ZN(n_1_232));
   AOI22_X1 i_1_400 (.A1(n_1_679), .A2(n_1_616), .B1(n_1_654), .B2(n_1_248), 
      .ZN(n_1_233));
   OAI221_X1 i_1_401 (.A(n_1_235), .B1(n_1_664), .B2(n_1_516), .C1(n_1_724), 
      .C2(n_1_629), .ZN(n_1_234));
   INV_X1 i_1_402 (.A(n_1_236), .ZN(n_1_235));
   OAI22_X1 i_1_403 (.A1(n_1_704), .A2(n_1_596), .B1(n_1_713), .B2(n_1_605), 
      .ZN(n_1_236));
   OR4_X1 i_1_404 (.A1(n_1_244), .A2(n_1_243), .A3(n_1_245), .A4(n_1_237), 
      .ZN(n_237));
   OR4_X1 i_1_405 (.A1(n_1_239), .A2(n_1_238), .A3(n_1_240), .A4(n_1_242), 
      .ZN(n_1_237));
   OAI22_X1 i_1_406 (.A1(n_1_534), .A2(n_1_516), .B1(n_1_656), .B2(n_1_531), 
      .ZN(n_1_238));
   OAI22_X1 i_1_407 (.A1(n_1_578), .A2(n_1_504), .B1(n_1_701), .B2(n_1_566), 
      .ZN(n_1_239));
   OAI221_X1 i_1_408 (.A(n_1_241), .B1(n_1_704), .B2(n_1_538), .C1(n_1_617), 
      .C2(n_1_575), .ZN(n_1_240));
   AOI22_X1 i_1_409 (.A1(n_1_725), .A2(n_1_551), .B1(n_1_648), .B2(n_1_548), 
      .ZN(n_1_241));
   OAI21_X1 i_1_410 (.A(n_1_694), .B1(n_1_727), .B2(n_1_721), .ZN(n_1_242));
   OAI22_X1 i_1_411 (.A1(n_1_707), .A2(n_1_560), .B1(n_1_645), .B2(n_1_541), 
      .ZN(n_1_243));
   OAI22_X1 i_1_412 (.A1(n_1_713), .A2(n_1_556), .B1(n_1_621), .B2(n_1_584), 
      .ZN(n_1_244));
   OAI221_X1 i_1_413 (.A(n_1_246), .B1(n_1_692), .B2(n_1_572), .C1(n_1_563), 
      .C2(n_1_247), .ZN(n_1_245));
   AOI22_X1 i_1_414 (.A1(n_1_662), .A2(n_1_582), .B1(n_1_554), .B2(n_1_487), 
      .ZN(n_1_246));
   INV_X1 i_1_415 (.A(n_1_248), .ZN(n_1_247));
   NOR3_X1 i_1_416 (.A1(counter[2]), .A2(n_1_717), .A3(n_1_722), .ZN(n_1_248));
   OR4_X1 i_1_417 (.A1(n_1_257), .A2(n_1_254), .A3(n_1_249), .A4(n_1_592), 
      .ZN(n_238));
   OR4_X1 i_1_418 (.A1(n_1_253), .A2(n_1_252), .A3(n_1_251), .A4(n_1_250), 
      .ZN(n_1_249));
   OAI22_X1 i_1_419 (.A1(n_1_701), .A2(n_1_596), .B1(n_1_664), .B2(n_1_504), 
      .ZN(n_1_250));
   OAI22_X1 i_1_420 (.A1(n_1_724), .A2(n_1_670), .B1(n_1_647), .B2(n_1_625), 
      .ZN(n_1_251));
   OAI22_X1 i_1_421 (.A1(n_1_678), .A2(n_1_656), .B1(n_1_707), .B2(n_1_618), 
      .ZN(n_1_252));
   NOR2_X1 i_1_422 (.A1(n_1_649), .A2(n_1_516), .ZN(n_1_253));
   OAI221_X1 i_1_423 (.A(n_1_255), .B1(n_1_617), .B2(n_1_600), .C1(n_1_674), 
      .C2(n_1_621), .ZN(n_1_254));
   INV_X1 i_1_424 (.A(n_1_256), .ZN(n_1_255));
   OAI22_X1 i_1_425 (.A1(n_1_704), .A2(n_1_609), .B1(n_1_713), .B2(n_1_637), 
      .ZN(n_1_256));
   OAI221_X1 i_1_426 (.A(n_1_258), .B1(n_1_605), .B2(n_1_486), .C1(n_1_661), 
      .C2(n_1_629), .ZN(n_1_257));
   INV_X1 i_1_427 (.A(n_1_259), .ZN(n_1_258));
   OAI22_X1 i_1_428 (.A1(n_1_684), .A2(n_1_645), .B1(n_1_692), .B2(n_1_653), 
      .ZN(n_1_259));
   OR4_X1 i_1_429 (.A1(n_1_262), .A2(n_1_260), .A3(n_1_264), .A4(n_1_592), 
      .ZN(n_239));
   OAI221_X1 i_1_430 (.A(n_1_261), .B1(n_1_692), .B2(n_1_563), .C1(n_1_701), 
      .C2(n_1_538), .ZN(n_1_260));
   AOI22_X1 i_1_431 (.A1(n_1_648), .A2(n_1_542), .B1(n_1_622), .B2(n_1_532), 
      .ZN(n_1_261));
   OAI221_X1 i_1_432 (.A(n_1_263), .B1(n_1_645), .B2(n_1_581), .C1(n_1_556), 
      .C2(n_1_486), .ZN(n_1_262));
   AOI22_X1 i_1_433 (.A1(n_1_712), .A2(n_1_561), .B1(n_1_708), .B2(n_1_573), 
      .ZN(n_1_263));
   OR4_X1 i_1_434 (.A1(n_1_268), .A2(n_1_267), .A3(n_1_266), .A4(n_1_265), 
      .ZN(n_1_264));
   OAI22_X1 i_1_435 (.A1(n_1_704), .A2(n_1_553), .B1(n_1_661), .B2(n_1_550), 
      .ZN(n_1_265));
   OAI22_X1 i_1_436 (.A1(n_1_547), .A2(n_1_516), .B1(n_1_640), .B2(n_1_584), 
      .ZN(n_1_266));
   OAI22_X1 i_1_437 (.A1(n_1_656), .A2(n_1_575), .B1(n_1_617), .B2(n_1_578), 
      .ZN(n_1_267));
   OAI22_X1 i_1_438 (.A1(n_1_724), .A2(n_1_566), .B1(n_1_534), .B2(n_1_504), 
      .ZN(n_1_268));
   OR4_X1 i_1_439 (.A1(n_1_276), .A2(n_1_274), .A3(n_1_269), .A4(n_1_591), 
      .ZN(n_240));
   OR4_X1 i_1_440 (.A1(n_1_273), .A2(n_1_272), .A3(n_1_271), .A4(n_1_270), 
      .ZN(n_1_269));
   OAI22_X1 i_1_441 (.A1(n_1_674), .A2(n_1_640), .B1(n_1_701), .B2(n_1_609), 
      .ZN(n_1_270));
   OAI22_X1 i_1_442 (.A1(n_1_678), .A2(n_1_621), .B1(n_1_704), .B2(n_1_605), 
      .ZN(n_1_271));
   OAI22_X1 i_1_443 (.A1(n_1_649), .A2(n_1_504), .B1(n_1_656), .B2(n_1_600), 
      .ZN(n_1_272));
   NOR2_X1 i_1_444 (.A1(n_1_645), .A2(n_1_629), .ZN(n_1_273));
   OAI221_X1 i_1_445 (.A(n_1_275), .B1(n_1_664), .B2(n_1_617), .C1(n_1_713), 
      .C2(n_1_618), .ZN(n_1_274));
   AOI22_X1 i_1_446 (.A1(n_1_725), .A2(n_1_597), .B1(n_1_638), .B2(n_1_487), 
      .ZN(n_1_275));
   OAI221_X1 i_1_447 (.A(n_1_277), .B1(n_1_670), .B2(n_1_661), .C1(n_1_625), 
      .C2(n_1_516), .ZN(n_1_276));
   AOI22_X1 i_1_448 (.A1(n_1_685), .A2(n_1_648), .B1(n_1_708), .B2(n_1_654), 
      .ZN(n_1_277));
   OR3_X1 i_1_449 (.A1(n_1_285), .A2(n_1_278), .A3(n_1_298), .ZN(n_241));
   OR4_X1 i_1_450 (.A1(n_1_280), .A2(n_1_279), .A3(n_1_281), .A4(n_1_284), 
      .ZN(n_1_278));
   OAI22_X1 i_1_451 (.A1(n_1_713), .A2(n_1_572), .B1(n_1_661), .B2(n_1_566), 
      .ZN(n_1_279));
   OAI22_X1 i_1_452 (.A1(n_1_541), .A2(n_1_516), .B1(n_1_707), .B2(n_1_563), 
      .ZN(n_1_280));
   OAI221_X1 i_1_453 (.A(n_1_282), .B1(n_1_656), .B2(n_1_578), .C1(n_1_701), 
      .C2(n_1_553), .ZN(n_1_281));
   INV_X1 i_1_454 (.A(n_1_283), .ZN(n_1_282));
   OAI22_X1 i_1_455 (.A1(n_1_560), .A2(n_1_486), .B1(n_1_640), .B2(n_1_531), 
      .ZN(n_1_283));
   OAI222_X1 i_1_456 (.A1(n_1_724), .A2(n_1_538), .B1(n_1_617), .B2(n_1_534), 
      .C1(n_1_547), .C2(n_1_504), .ZN(n_1_284));
   OAI211_X1 i_1_457 (.A(n_1_698), .B(n_1_286), .C1(n_1_608), .C2(n_1_584), 
      .ZN(n_1_285));
   AOI221_X1 i_1_458 (.A(n_1_287), .B1(n_1_622), .B2(n_1_576), .C1(n_1_648), 
      .C2(n_1_582), .ZN(n_1_286));
   OAI22_X1 i_1_459 (.A1(n_1_704), .A2(n_1_556), .B1(n_1_645), .B2(n_1_550), 
      .ZN(n_1_287));
   OR3_X1 i_1_460 (.A1(n_1_295), .A2(n_1_288), .A3(n_1_298), .ZN(n_242));
   OR4_X1 i_1_461 (.A1(n_1_290), .A2(n_1_289), .A3(n_1_291), .A4(n_1_294), 
      .ZN(n_1_288));
   OAI22_X1 i_1_462 (.A1(n_1_618), .A2(n_1_486), .B1(n_1_704), .B2(n_1_637), 
      .ZN(n_1_289));
   OAI22_X1 i_1_463 (.A1(n_1_684), .A2(n_1_516), .B1(n_1_701), .B2(n_1_605), 
      .ZN(n_1_290));
   OAI221_X1 i_1_464 (.A(n_1_292), .B1(n_1_664), .B2(n_1_656), .C1(n_1_674), 
      .C2(n_1_608), .ZN(n_1_291));
   INV_X1 i_1_465 (.A(n_1_293), .ZN(n_1_292));
   OAI22_X1 i_1_466 (.A1(n_1_678), .A2(n_1_640), .B1(n_1_670), .B2(n_1_645), 
      .ZN(n_1_293));
   OAI222_X1 i_1_467 (.A1(n_1_661), .A2(n_1_596), .B1(n_1_625), .B2(n_1_504), 
      .C1(n_1_724), .C2(n_1_609), .ZN(n_1_294));
   OR4_X1 i_1_468 (.A1(n_1_706), .A2(n_1_699), .A3(n_1_297), .A4(n_1_296), 
      .ZN(n_1_295));
   OAI22_X1 i_1_469 (.A1(n_1_713), .A2(n_1_653), .B1(n_1_649), .B2(n_1_617), 
      .ZN(n_1_296));
   OAI22_X1 i_1_470 (.A1(n_1_647), .A2(n_1_629), .B1(n_1_621), .B2(n_1_600), 
      .ZN(n_1_297));
   OR2_X1 i_1_471 (.A1(n_1_695), .A2(n_1_393), .ZN(n_1_298));
   OR4_X1 i_1_472 (.A1(n_1_693), .A2(n_1_306), .A3(n_1_299), .A4(n_1_392), 
      .ZN(n_243));
   OR4_X1 i_1_473 (.A1(n_1_301), .A2(n_1_300), .A3(n_1_302), .A4(n_1_304), 
      .ZN(n_1_299));
   OAI22_X1 i_1_474 (.A1(n_1_640), .A2(n_1_575), .B1(n_1_647), .B2(n_1_550), 
      .ZN(n_1_300));
   OAI22_X1 i_1_475 (.A1(n_1_656), .A2(n_1_534), .B1(n_1_701), .B2(n_1_556), 
      .ZN(n_1_301));
   OAI221_X1 i_1_476 (.A(n_1_303), .B1(n_1_621), .B2(n_1_578), .C1(n_1_704), 
      .C2(n_1_560), .ZN(n_1_302));
   AOI22_X1 i_1_477 (.A1(n_1_582), .A2(n_1_517), .B1(n_1_573), .B2(n_1_487), 
      .ZN(n_1_303));
   OAI221_X1 i_1_478 (.A(n_1_305), .B1(n_1_661), .B2(n_1_538), .C1(n_1_724), 
      .C2(n_1_553), .ZN(n_1_304));
   AOI22_X1 i_1_479 (.A1(n_1_542), .A2(n_1_505), .B1(n_1_712), .B2(n_1_564), 
      .ZN(n_1_305));
   OAI221_X1 i_1_480 (.A(n_1_307), .B1(n_1_617), .B2(n_1_547), .C1(n_1_612), 
      .C2(n_1_584), .ZN(n_1_306));
   INV_X1 i_1_481 (.A(n_1_308), .ZN(n_1_307));
   OAI22_X1 i_1_482 (.A1(n_1_608), .A2(n_1_531), .B1(n_1_645), .B2(n_1_566), 
      .ZN(n_1_308));
   OR4_X1 i_1_483 (.A1(n_1_693), .A2(n_1_317), .A3(n_1_309), .A4(n_1_392), 
      .ZN(n_244));
   OR4_X1 i_1_484 (.A1(n_1_311), .A2(n_1_310), .A3(n_1_312), .A4(n_1_315), 
      .ZN(n_1_309));
   OAI22_X1 i_1_485 (.A1(n_1_653), .A2(n_1_486), .B1(n_1_674), .B2(n_1_612), 
      .ZN(n_1_310));
   OAI22_X1 i_1_486 (.A1(n_1_645), .A2(n_1_596), .B1(n_1_670), .B2(n_1_647), 
      .ZN(n_1_311));
   OAI221_X1 i_1_487 (.A(n_1_313), .B1(n_1_684), .B2(n_1_504), .C1(n_1_701), 
      .C2(n_1_637), .ZN(n_1_312));
   INV_X1 i_1_488 (.A(n_1_314), .ZN(n_1_313));
   OAI22_X1 i_1_489 (.A1(n_1_678), .A2(n_1_608), .B1(n_1_704), .B2(n_1_618), 
      .ZN(n_1_314));
   OAI221_X1 i_1_490 (.A(n_1_316), .B1(n_1_724), .B2(n_1_605), .C1(n_1_625), 
      .C2(n_1_617), .ZN(n_1_315));
   AOI22_X1 i_1_491 (.A1(n_1_662), .A2(n_1_610), .B1(n_1_630), .B2(n_1_517), 
      .ZN(n_1_316));
   OAI221_X1 i_1_492 (.A(n_1_318), .B1(n_1_640), .B2(n_1_600), .C1(n_1_664), 
      .C2(n_1_621), .ZN(n_1_317));
   INV_X1 i_1_493 (.A(n_1_319), .ZN(n_1_318));
   OAI21_X1 i_1_494 (.A(n_1_710), .B1(n_1_656), .B2(n_1_649), .ZN(n_1_319));
   OR4_X1 i_1_495 (.A1(n_1_705), .A2(n_1_327), .A3(n_1_320), .A4(n_1_591), 
      .ZN(n_245));
   OR4_X1 i_1_496 (.A1(n_1_324), .A2(n_1_323), .A3(n_1_321), .A4(n_1_325), 
      .ZN(n_1_320));
   OAI221_X1 i_1_497 (.A(n_1_322), .B1(n_1_640), .B2(n_1_578), .C1(n_1_704), 
      .C2(n_1_572), .ZN(n_1_321));
   AOI22_X1 i_1_498 (.A1(n_1_646), .A2(n_1_539), .B1(n_1_648), .B2(n_1_567), 
      .ZN(n_1_322));
   OAI22_X1 i_1_499 (.A1(n_1_612), .A2(n_1_531), .B1(n_1_621), .B2(n_1_534), 
      .ZN(n_1_323));
   OAI22_X1 i_1_500 (.A1(n_1_617), .A2(n_1_541), .B1(n_1_701), .B2(n_1_560), 
      .ZN(n_1_324));
   OAI221_X1 i_1_501 (.A(n_1_326), .B1(n_1_550), .B2(n_1_516), .C1(n_1_656), 
      .C2(n_1_547), .ZN(n_1_325));
   AOI22_X1 i_1_502 (.A1(n_1_662), .A2(n_1_554), .B1(n_1_564), .B2(n_1_487), 
      .ZN(n_1_326));
   OAI221_X1 i_1_503 (.A(n_1_328), .B1(n_1_581), .B2(n_1_504), .C1(n_1_724), 
      .C2(n_1_556), .ZN(n_1_327));
   INV_X1 i_1_504 (.A(n_1_329), .ZN(n_1_328));
   OAI22_X1 i_1_505 (.A1(n_1_608), .A2(n_1_575), .B1(n_1_599), .B2(n_1_584), 
      .ZN(n_1_329));
   OR4_X1 i_1_506 (.A1(n_1_337), .A2(n_1_335), .A3(n_1_330), .A4(n_1_588), 
      .ZN(n_246));
   OR4_X1 i_1_507 (.A1(n_1_334), .A2(n_1_333), .A3(n_1_332), .A4(n_1_331), 
      .ZN(n_1_330));
   OAI22_X1 i_1_508 (.A1(n_1_704), .A2(n_1_653), .B1(n_1_647), .B2(n_1_596), 
      .ZN(n_1_331));
   OAI22_X1 i_1_509 (.A1(n_1_678), .A2(n_1_612), .B1(n_1_608), .B2(n_1_600), 
      .ZN(n_1_332));
   OAI22_X1 i_1_510 (.A1(n_1_701), .A2(n_1_618), .B1(n_1_664), .B2(n_1_640), 
      .ZN(n_1_333));
   NOR2_X1 i_1_511 (.A1(n_1_674), .A2(n_1_599), .ZN(n_1_334));
   OAI221_X1 i_1_512 (.A(n_1_336), .B1(n_1_656), .B2(n_1_625), .C1(n_1_670), 
      .C2(n_1_516), .ZN(n_1_335));
   AOI22_X1 i_1_513 (.A1(n_1_725), .A2(n_1_638), .B1(n_1_650), .B2(n_1_622), 
      .ZN(n_1_336));
   OAI221_X1 i_1_514 (.A(n_1_338), .B1(n_1_629), .B2(n_1_504), .C1(n_1_684), 
      .C2(n_1_617), .ZN(n_1_337));
   AOI22_X1 i_1_515 (.A1(n_1_662), .A2(n_1_606), .B1(n_1_646), .B2(n_1_610), 
      .ZN(n_1_338));
   OR4_X1 i_1_516 (.A1(n_1_342), .A2(n_1_339), .A3(n_1_344), .A4(n_1_588), 
      .ZN(n_247));
   OAI221_X1 i_1_517 (.A(n_1_340), .B1(n_1_612), .B2(n_1_575), .C1(n_1_661), 
      .C2(n_1_556), .ZN(n_1_339));
   INV_X1 i_1_518 (.A(n_1_341), .ZN(n_1_340));
   OAI22_X1 i_1_519 (.A1(n_1_701), .A2(n_1_572), .B1(n_1_704), .B2(n_1_563), 
      .ZN(n_1_341));
   OAI221_X1 i_1_520 (.A(n_1_343), .B1(n_1_608), .B2(n_1_578), .C1(n_1_550), 
      .C2(n_1_504), .ZN(n_1_342));
   AOI22_X1 i_1_521 (.A1(n_1_646), .A2(n_1_554), .B1(n_1_567), .B2(n_1_517), 
      .ZN(n_1_343));
   OR4_X1 i_1_522 (.A1(n_1_348), .A2(n_1_347), .A3(n_1_346), .A4(n_1_345), 
      .ZN(n_1_344));
   OAI22_X1 i_1_523 (.A1(n_1_724), .A2(n_1_560), .B1(n_1_621), .B2(n_1_547), 
      .ZN(n_1_345));
   OAI22_X1 i_1_524 (.A1(n_1_599), .A2(n_1_531), .B1(n_1_673), .B2(n_1_584), 
      .ZN(n_1_346));
   OAI22_X1 i_1_525 (.A1(n_1_656), .A2(n_1_541), .B1(n_1_617), .B2(n_1_581), 
      .ZN(n_1_347));
   OAI22_X1 i_1_526 (.A1(n_1_640), .A2(n_1_534), .B1(n_1_647), .B2(n_1_538), 
      .ZN(n_1_348));
   OR4_X1 i_1_527 (.A1(n_1_356), .A2(n_1_353), .A3(n_1_349), .A4(n_1_370), 
      .ZN(n_248));
   OR4_X1 i_1_528 (.A1(n_1_351), .A2(n_1_350), .A3(n_1_352), .A4(n_1_593), 
      .ZN(n_1_349));
   OAI22_X1 i_1_529 (.A1(n_1_629), .A2(n_1_617), .B1(n_1_625), .B2(n_1_621), 
      .ZN(n_1_350));
   OAI22_X1 i_1_530 (.A1(n_1_596), .A2(n_1_516), .B1(n_1_670), .B2(n_1_504), 
      .ZN(n_1_351));
   OAI222_X1 i_1_531 (.A1(n_1_612), .A2(n_1_600), .B1(n_1_674), .B2(n_1_673), 
      .C1(n_1_647), .C2(n_1_609), .ZN(n_1_352));
   OAI221_X1 i_1_532 (.A(n_1_354), .B1(n_1_684), .B2(n_1_656), .C1(n_1_664), 
      .C2(n_1_608), .ZN(n_1_353));
   INV_X1 i_1_533 (.A(n_1_355), .ZN(n_1_354));
   OAI22_X1 i_1_534 (.A1(n_1_649), .A2(n_1_640), .B1(n_1_645), .B2(n_1_605), 
      .ZN(n_1_355));
   OAI221_X1 i_1_535 (.A(n_1_357), .B1(n_1_661), .B2(n_1_637), .C1(n_1_724), 
      .C2(n_1_618), .ZN(n_1_356));
   INV_X1 i_1_536 (.A(n_1_358), .ZN(n_1_357));
   OAI22_X1 i_1_537 (.A1(n_1_701), .A2(n_1_653), .B1(n_1_678), .B2(n_1_599), 
      .ZN(n_1_358));
   OR4_X1 i_1_538 (.A1(n_1_367), .A2(n_1_364), .A3(n_1_359), .A4(n_1_370), 
      .ZN(n_249));
   OR4_X1 i_1_539 (.A1(n_1_361), .A2(n_1_360), .A3(n_1_362), .A4(n_1_593), 
      .ZN(n_1_359));
   OAI22_X1 i_1_540 (.A1(n_1_599), .A2(n_1_575), .B1(n_1_612), .B2(n_1_578), 
      .ZN(n_1_360));
   OAI22_X1 i_1_541 (.A1(n_1_538), .A2(n_1_516), .B1(n_1_640), .B2(n_1_547), 
      .ZN(n_1_361));
   OAI221_X1 i_1_542 (.A(n_1_363), .B1(n_1_701), .B2(n_1_563), .C1(n_1_656), 
      .C2(n_1_581), .ZN(n_1_362));
   AOI22_X1 i_1_543 (.A1(n_1_662), .A2(n_1_561), .B1(n_1_646), .B2(n_1_557), 
      .ZN(n_1_363));
   OAI221_X1 i_1_544 (.A(n_1_365), .B1(n_1_724), .B2(n_1_572), .C1(n_1_608), 
      .C2(n_1_534), .ZN(n_1_364));
   INV_X1 i_1_545 (.A(n_1_366), .ZN(n_1_365));
   OAI22_X1 i_1_546 (.A1(n_1_647), .A2(n_1_553), .B1(n_1_632), .B2(n_1_584), 
      .ZN(n_1_366));
   OAI221_X1 i_1_547 (.A(n_1_368), .B1(n_1_617), .B2(n_1_550), .C1(n_1_621), 
      .C2(n_1_541), .ZN(n_1_367));
   INV_X1 i_1_548 (.A(n_1_369), .ZN(n_1_368));
   OAI22_X1 i_1_549 (.A1(n_1_566), .A2(n_1_504), .B1(n_1_673), .B2(n_1_531), 
      .ZN(n_1_369));
   OR3_X1 i_1_550 (.A1(n_1_703), .A2(n_1_690), .A3(n_1_589), .ZN(n_1_370));
   NAND3_X1 i_1_551 (.A1(n_1_689), .A2(n_1_371), .A3(n_1_376), .ZN(n_250));
   NOR4_X1 i_1_552 (.A1(n_1_375), .A2(n_1_374), .A3(n_1_373), .A4(n_1_372), 
      .ZN(n_1_371));
   OAI22_X1 i_1_553 (.A1(n_1_674), .A2(n_1_632), .B1(n_1_656), .B2(n_1_629), 
      .ZN(n_1_372));
   OAI22_X1 i_1_554 (.A1(n_1_670), .A2(n_1_617), .B1(n_1_724), .B2(n_1_653), 
      .ZN(n_1_373));
   OAI22_X1 i_1_555 (.A1(n_1_678), .A2(n_1_673), .B1(n_1_596), .B2(n_1_504), 
      .ZN(n_1_374));
   OAI22_X1 i_1_556 (.A1(n_1_640), .A2(n_1_625), .B1(n_1_609), .B2(n_1_516), 
      .ZN(n_1_375));
   NOR4_X1 i_1_557 (.A1(n_1_378), .A2(n_1_377), .A3(n_1_379), .A4(n_1_719), 
      .ZN(n_1_376));
   OAI22_X1 i_1_558 (.A1(n_1_684), .A2(n_1_621), .B1(n_1_649), .B2(n_1_608), 
      .ZN(n_1_377));
   OAI22_X1 i_1_559 (.A1(n_1_600), .A2(n_1_599), .B1(n_1_647), .B2(n_1_605), 
      .ZN(n_1_378));
   OAI222_X1 i_1_560 (.A1(n_1_664), .A2(n_1_612), .B1(n_1_645), .B2(n_1_637), 
      .C1(n_1_661), .C2(n_1_618), .ZN(n_1_379));
   OR3_X1 i_1_561 (.A1(n_1_383), .A2(n_1_380), .A3(n_1_392), .ZN(n_251));
   OR3_X1 i_1_562 (.A1(n_1_693), .A2(n_1_381), .A3(n_1_404), .ZN(n_1_380));
   OAI221_X1 i_1_563 (.A(n_1_382), .B1(n_1_640), .B2(n_1_541), .C1(n_1_687), 
      .C2(n_1_584), .ZN(n_1_381));
   AOI22_X1 i_1_564 (.A1(n_1_662), .A2(n_1_573), .B1(n_1_646), .B2(n_1_561), 
      .ZN(n_1_382));
   OR4_X1 i_1_565 (.A1(n_1_385), .A2(n_1_384), .A3(n_1_386), .A4(n_1_389), 
      .ZN(n_1_383));
   OAI22_X1 i_1_566 (.A1(n_1_599), .A2(n_1_578), .B1(n_1_553), .B2(n_1_516), 
      .ZN(n_1_384));
   OAI22_X1 i_1_567 (.A1(n_1_647), .A2(n_1_556), .B1(n_1_632), .B2(n_1_531), 
      .ZN(n_1_385));
   OAI221_X1 i_1_568 (.A(n_1_387), .B1(n_1_621), .B2(n_1_581), .C1(n_1_608), 
      .C2(n_1_547), .ZN(n_1_386));
   INV_X1 i_1_569 (.A(n_1_388), .ZN(n_1_387));
   OAI22_X1 i_1_570 (.A1(n_1_656), .A2(n_1_550), .B1(n_1_673), .B2(n_1_575), 
      .ZN(n_1_388));
   OAI221_X1 i_1_571 (.A(n_1_390), .B1(n_1_538), .B2(n_1_504), .C1(n_1_617), 
      .C2(n_1_566), .ZN(n_1_389));
   INV_X1 i_1_572 (.A(n_1_391), .ZN(n_1_390));
   OAI22_X1 i_1_573 (.A1(n_1_612), .A2(n_1_534), .B1(n_1_724), .B2(n_1_563), 
      .ZN(n_1_391));
   OR2_X1 i_1_574 (.A1(n_1_706), .A2(n_1_393), .ZN(n_1_392));
   OR2_X1 i_1_575 (.A1(n_1_691), .A2(n_1_593), .ZN(n_1_393));
   OR4_X1 i_1_576 (.A1(n_1_690), .A2(n_1_405), .A3(n_1_593), .A4(n_1_394), 
      .ZN(n_252));
   OR4_X1 i_1_577 (.A1(n_1_398), .A2(n_1_395), .A3(n_1_401), .A4(n_1_404), 
      .ZN(n_1_394));
   OAI221_X1 i_1_578 (.A(n_1_396), .B1(n_1_684), .B2(n_1_640), .C1(n_1_605), 
      .C2(n_1_516), .ZN(n_1_395));
   INV_X1 i_1_579 (.A(n_1_397), .ZN(n_1_396));
   OAI22_X1 i_1_580 (.A1(n_1_687), .A2(n_1_674), .B1(n_1_670), .B2(n_1_656), 
      .ZN(n_1_397));
   OAI221_X1 i_1_581 (.A(n_1_399), .B1(n_1_629), .B2(n_1_621), .C1(n_1_617), 
      .C2(n_1_596), .ZN(n_1_398));
   INV_X1 i_1_582 (.A(n_1_400), .ZN(n_1_399));
   OAI22_X1 i_1_583 (.A1(n_1_609), .A2(n_1_504), .B1(n_1_673), .B2(n_1_600), 
      .ZN(n_1_400));
   OR4_X1 i_1_584 (.A1(n_1_723), .A2(n_1_706), .A3(n_1_403), .A4(n_1_402), 
      .ZN(n_1_401));
   OAI22_X1 i_1_585 (.A1(n_1_645), .A2(n_1_618), .B1(n_1_664), .B2(n_1_599), 
      .ZN(n_1_402));
   OAI22_X1 i_1_586 (.A1(n_1_647), .A2(n_1_637), .B1(n_1_649), .B2(n_1_612), 
      .ZN(n_1_403));
   OR3_X1 i_1_587 (.A1(n_1_711), .A2(n_1_938), .A3(n_1_590), .ZN(n_1_404));
   OAI222_X1 i_1_588 (.A1(n_1_661), .A2(n_1_653), .B1(n_1_678), .B2(n_1_632), 
      .C1(n_1_625), .C2(n_1_608), .ZN(n_1_405));
   OR4_X1 i_1_589 (.A1(n_1_408), .A2(n_1_406), .A3(n_1_411), .A4(n_1_688), 
      .ZN(n_253));
   OAI221_X1 i_1_590 (.A(n_1_407), .B1(n_1_599), .B2(n_1_534), .C1(n_1_640), 
      .C2(n_1_581), .ZN(n_1_406));
   AOI22_X1 i_1_591 (.A1(n_1_633), .A2(n_1_576), .B1(n_1_646), .B2(n_1_573), 
      .ZN(n_1_407));
   OAI221_X1 i_1_592 (.A(n_1_409), .B1(n_1_612), .B2(n_1_547), .C1(n_1_617), 
      .C2(n_1_538), .ZN(n_1_408));
   INV_X1 i_1_593 (.A(n_1_410), .ZN(n_1_409));
   OAI22_X1 i_1_594 (.A1(n_1_608), .A2(n_1_541), .B1(n_1_656), .B2(n_1_566), 
      .ZN(n_1_410));
   OR4_X1 i_1_595 (.A1(n_1_415), .A2(n_1_414), .A3(n_1_413), .A4(n_1_412), 
      .ZN(n_1_411));
   OAI22_X1 i_1_596 (.A1(n_1_673), .A2(n_1_578), .B1(n_1_553), .B2(n_1_504), 
      .ZN(n_1_412));
   OAI22_X1 i_1_597 (.A1(n_1_687), .A2(n_1_531), .B1(n_1_628), .B2(n_1_584), 
      .ZN(n_1_413));
   OAI22_X1 i_1_598 (.A1(n_1_621), .A2(n_1_550), .B1(n_1_647), .B2(n_1_560), 
      .ZN(n_1_414));
   OAI22_X1 i_1_599 (.A1(n_1_661), .A2(n_1_563), .B1(n_1_556), .B2(n_1_516), 
      .ZN(n_1_415));
   OR3_X1 i_1_600 (.A1(n_1_423), .A2(n_1_416), .A3(n_1_591), .ZN(n_254));
   OR4_X1 i_1_601 (.A1(n_1_420), .A2(n_1_418), .A3(n_1_700), .A4(n_1_417), 
      .ZN(n_1_416));
   OAI222_X1 i_1_602 (.A1(n_1_637), .A2(n_1_516), .B1(n_1_687), .B2(n_1_678), 
      .C1(n_1_684), .C2(n_1_608), .ZN(n_1_417));
   OAI221_X1 i_1_603 (.A(n_1_419), .B1(n_1_656), .B2(n_1_596), .C1(n_1_605), 
      .C2(n_1_504), .ZN(n_1_418));
   AOI22_X1 i_1_604 (.A1(n_1_616), .A2(n_1_610), .B1(n_1_633), .B2(n_1_601), 
      .ZN(n_1_419));
   OAI221_X1 i_1_605 (.A(n_1_421), .B1(n_1_647), .B2(n_1_618), .C1(n_1_625), 
      .C2(n_1_612), .ZN(n_1_420));
   INV_X1 i_1_606 (.A(n_1_422), .ZN(n_1_421));
   OAI22_X1 i_1_607 (.A1(n_1_653), .A2(n_1_645), .B1(n_1_649), .B2(n_1_599), 
      .ZN(n_1_422));
   OR4_X1 i_1_608 (.A1(n_1_425), .A2(n_1_424), .A3(n_1_590), .A4(n_1_587), 
      .ZN(n_1_423));
   OAI22_X1 i_1_609 (.A1(n_1_640), .A2(n_1_629), .B1(n_1_674), .B2(n_1_628), 
      .ZN(n_1_424));
   OAI22_X1 i_1_610 (.A1(n_1_670), .A2(n_1_621), .B1(n_1_673), .B2(n_1_664), 
      .ZN(n_1_425));
   OR4_X1 i_1_611 (.A1(n_1_429), .A2(n_1_426), .A3(n_1_432), .A4(n_1_585), 
      .ZN(n_255));
   OAI221_X1 i_1_612 (.A(n_1_427), .B1(n_1_647), .B2(n_1_572), .C1(n_1_640), 
      .C2(n_1_550), .ZN(n_1_426));
   INV_X1 i_1_613 (.A(n_1_428), .ZN(n_1_427));
   OAI22_X1 i_1_614 (.A1(n_1_687), .A2(n_1_575), .B1(n_1_656), .B2(n_1_538), 
      .ZN(n_1_428));
   OAI221_X1 i_1_615 (.A(n_1_430), .B1(n_1_608), .B2(n_1_581), .C1(n_1_560), 
      .C2(n_1_516), .ZN(n_1_429));
   INV_X1 i_1_616 (.A(n_1_431), .ZN(n_1_430));
   OAI22_X1 i_1_617 (.A1(n_1_599), .A2(n_1_547), .B1(n_1_612), .B2(n_1_541), 
      .ZN(n_1_431));
   OR4_X1 i_1_618 (.A1(n_1_436), .A2(n_1_435), .A3(n_1_434), .A4(n_1_433), 
      .ZN(n_1_432));
   OAI22_X1 i_1_619 (.A1(n_1_628), .A2(n_1_531), .B1(n_1_556), .B2(n_1_504), 
      .ZN(n_1_433));
   OAI22_X1 i_1_620 (.A1(n_1_617), .A2(n_1_553), .B1(n_1_652), .B2(n_1_584), 
      .ZN(n_1_434));
   OAI22_X1 i_1_621 (.A1(n_1_632), .A2(n_1_578), .B1(n_1_645), .B2(n_1_563), 
      .ZN(n_1_435));
   OAI22_X1 i_1_622 (.A1(n_1_621), .A2(n_1_566), .B1(n_1_673), .B2(n_1_534), 
      .ZN(n_1_436));
   OR4_X1 i_1_623 (.A1(n_1_705), .A2(n_1_446), .A3(n_1_437), .A4(n_1_591), 
      .ZN(n_256));
   OR4_X1 i_1_624 (.A1(n_1_443), .A2(n_1_441), .A3(n_1_586), .A4(n_1_438), 
      .ZN(n_1_437));
   OAI221_X1 i_1_625 (.A(n_1_439), .B1(n_1_629), .B2(n_1_608), .C1(n_1_670), 
      .C2(n_1_640), .ZN(n_1_438));
   INV_X1 i_1_626 (.A(n_1_440), .ZN(n_1_439));
   OAI22_X1 i_1_627 (.A1(n_1_673), .A2(n_1_649), .B1(n_1_684), .B2(n_1_612), 
      .ZN(n_1_440));
   OAI221_X1 i_1_628 (.A(n_1_442), .B1(n_1_621), .B2(n_1_596), .C1(n_1_674), 
      .C2(n_1_652), .ZN(n_1_441));
   AOI22_X1 i_1_629 (.A1(n_1_616), .A2(n_1_606), .B1(n_1_619), .B2(n_1_517), 
      .ZN(n_1_442));
   OAI221_X1 i_1_630 (.A(n_1_444), .B1(n_1_656), .B2(n_1_609), .C1(n_1_637), 
      .C2(n_1_504), .ZN(n_1_443));
   INV_X1 i_1_631 (.A(n_1_445), .ZN(n_1_444));
   OAI22_X1 i_1_632 (.A1(n_1_678), .A2(n_1_628), .B1(n_1_653), .B2(n_1_647), 
      .ZN(n_1_445));
   OAI221_X1 i_1_633 (.A(n_1_447), .B1(n_1_664), .B2(n_1_632), .C1(n_1_687), 
      .C2(n_1_600), .ZN(n_1_446));
   INV_X1 i_1_634 (.A(n_1_448), .ZN(n_1_447));
   OAI21_X1 i_1_635 (.A(n_1_455), .B1(n_1_625), .B2(n_1_599), .ZN(n_1_448));
   NAND3_X1 i_1_636 (.A1(n_1_488), .A2(n_1_449), .A3(n_1_459), .ZN(n_257));
   NOR4_X1 i_1_637 (.A1(n_1_451), .A2(n_1_450), .A3(n_1_452), .A4(n_1_456), 
      .ZN(n_1_449));
   OAI22_X1 i_1_638 (.A1(n_1_628), .A2(n_1_575), .B1(n_1_673), .B2(n_1_547), 
      .ZN(n_1_450));
   OAI22_X1 i_1_639 (.A1(n_1_621), .A2(n_1_538), .B1(n_1_647), .B2(n_1_563), 
      .ZN(n_1_451));
   OAI221_X1 i_1_640 (.A(n_1_453), .B1(n_1_656), .B2(n_1_553), .C1(n_1_640), 
      .C2(n_1_566), .ZN(n_1_452));
   INV_X1 i_1_641 (.A(n_1_454), .ZN(n_1_453));
   OAI21_X1 i_1_642 (.A(n_1_455), .B1(n_1_572), .B2(n_1_516), .ZN(n_1_454));
   OAI21_X1 i_1_643 (.A(n_1_729), .B1(n_1_646), .B2(n_1_487), .ZN(n_1_455));
   OAI221_X1 i_1_644 (.A(n_1_457), .B1(n_1_560), .B2(n_1_504), .C1(n_1_667), 
      .C2(n_1_584), .ZN(n_1_456));
   AOI221_X1 i_1_645 (.A(n_1_458), .B1(n_1_633), .B2(n_1_535), .C1(n_1_616), 
      .C2(n_1_557), .ZN(n_1_457));
   OAI22_X1 i_1_646 (.A1(n_1_612), .A2(n_1_581), .B1(n_1_687), .B2(n_1_578), 
      .ZN(n_1_458));
   NOR3_X1 i_1_647 (.A1(n_1_700), .A2(n_1_460), .A3(n_1_593), .ZN(n_1_459));
   OAI222_X1 i_1_648 (.A1(n_1_599), .A2(n_1_541), .B1(n_1_608), .B2(n_1_550), 
      .C1(n_1_652), .C2(n_1_531), .ZN(n_1_460));
   OR4_X1 i_1_649 (.A1(n_1_468), .A2(n_1_465), .A3(n_1_461), .A4(n_1_484), 
      .ZN(n_258));
   OR4_X1 i_1_650 (.A1(n_1_463), .A2(n_1_462), .A3(n_1_464), .A4(n_1_472), 
      .ZN(n_1_461));
   OAI22_X1 i_1_651 (.A1(n_1_674), .A2(n_1_667), .B1(n_1_618), .B2(n_1_504), 
      .ZN(n_1_462));
   OAI22_X1 i_1_652 (.A1(n_1_629), .A2(n_1_612), .B1(n_1_649), .B2(n_1_632), 
      .ZN(n_1_463));
   OAI222_X1 i_1_653 (.A1(n_1_628), .A2(n_1_600), .B1(n_1_640), .B2(n_1_596), 
      .C1(n_1_684), .C2(n_1_599), .ZN(n_1_464));
   OAI221_X1 i_1_654 (.A(n_1_466), .B1(n_1_656), .B2(n_1_605), .C1(n_1_621), 
      .C2(n_1_609), .ZN(n_1_465));
   INV_X1 i_1_655 (.A(n_1_467), .ZN(n_1_466));
   OAI22_X1 i_1_656 (.A1(n_1_687), .A2(n_1_664), .B1(n_1_637), .B2(n_1_617), 
      .ZN(n_1_467));
   OAI221_X1 i_1_657 (.A(n_1_469), .B1(n_1_673), .B2(n_1_625), .C1(n_1_670), 
      .C2(n_1_608), .ZN(n_1_468));
   INV_X1 i_1_658 (.A(n_1_470), .ZN(n_1_469));
   OAI22_X1 i_1_659 (.A1(n_1_678), .A2(n_1_652), .B1(n_1_653), .B2(n_1_516), 
      .ZN(n_1_470));
   OR4_X1 i_1_660 (.A1(n_1_481), .A2(n_1_478), .A3(n_1_471), .A4(n_1_484), 
      .ZN(n_259));
   OR4_X1 i_1_661 (.A1(n_1_474), .A2(n_1_473), .A3(n_1_475), .A4(n_1_472), 
      .ZN(n_1_471));
   OR2_X1 i_1_662 (.A1(n_1_700), .A2(n_1_593), .ZN(n_1_472));
   OAI22_X1 i_1_663 (.A1(n_1_656), .A2(n_1_556), .B1(n_1_563), .B2(n_1_516), 
      .ZN(n_1_473));
   OAI22_X1 i_1_664 (.A1(n_1_621), .A2(n_1_553), .B1(n_1_652), .B2(n_1_575), 
      .ZN(n_1_474));
   OAI221_X1 i_1_665 (.A(n_1_476), .B1(n_1_612), .B2(n_1_550), .C1(n_1_673), 
      .C2(n_1_541), .ZN(n_1_475));
   INV_X1 i_1_666 (.A(n_1_477), .ZN(n_1_476));
   OAI22_X1 i_1_667 (.A1(n_1_628), .A2(n_1_578), .B1(n_1_599), .B2(n_1_581), 
      .ZN(n_1_477));
   OAI221_X1 i_1_668 (.A(n_1_479), .B1(n_1_617), .B2(n_1_560), .C1(n_1_608), 
      .C2(n_1_566), .ZN(n_1_478));
   INV_X1 i_1_669 (.A(n_1_480), .ZN(n_1_479));
   OAI22_X1 i_1_670 (.A1(n_1_667), .A2(n_1_531), .B1(n_1_603), .B2(n_1_584), 
      .ZN(n_1_480));
   OAI221_X1 i_1_671 (.A(n_1_482), .B1(n_1_632), .B2(n_1_547), .C1(n_1_640), 
      .C2(n_1_538), .ZN(n_1_481));
   INV_X1 i_1_672 (.A(n_1_483), .ZN(n_1_482));
   OAI22_X1 i_1_673 (.A1(n_1_687), .A2(n_1_534), .B1(n_1_572), .B2(n_1_504), 
      .ZN(n_1_483));
   OAI21_X1 i_1_674 (.A(n_1_488), .B1(n_1_728), .B2(n_1_485), .ZN(n_1_484));
   NOR2_X1 i_1_675 (.A1(n_1_644), .A2(n_1_487), .ZN(n_1_485));
   INV_X1 i_1_676 (.A(n_1_487), .ZN(n_1_486));
   NOR2_X1 i_1_677 (.A1(n_1_722), .A2(n_1_716), .ZN(n_1_487));
   NOR2_X1 i_1_678 (.A1(n_1_690), .A2(n_1_587), .ZN(n_1_488));
   OR3_X1 i_1_679 (.A1(n_1_718), .A2(n_1_489), .A3(n_1_514), .ZN(n_260));
   OR4_X1 i_1_680 (.A1(n_1_496), .A2(n_1_494), .A3(n_1_493), .A4(n_1_490), 
      .ZN(n_1_489));
   OAI221_X1 i_1_681 (.A(n_1_491), .B1(n_1_687), .B2(n_1_649), .C1(n_1_670), 
      .C2(n_1_612), .ZN(n_1_490));
   INV_X1 i_1_682 (.A(n_1_492), .ZN(n_1_491));
   OAI22_X1 i_1_683 (.A1(n_1_678), .A2(n_1_667), .B1(n_1_640), .B2(n_1_609), 
      .ZN(n_1_492));
   OAI222_X1 i_1_684 (.A1(n_1_684), .A2(n_1_673), .B1(n_1_629), .B2(n_1_599), 
      .C1(n_1_608), .C2(n_1_596), .ZN(n_1_493));
   OAI221_X1 i_1_685 (.A(n_1_495), .B1(n_1_618), .B2(n_1_617), .C1(n_1_621), 
      .C2(n_1_605), .ZN(n_1_494));
   AOI22_X1 i_1_686 (.A1(n_1_654), .A2(n_1_505), .B1(n_1_633), .B2(n_1_626), 
      .ZN(n_1_495));
   OAI221_X1 i_1_687 (.A(n_1_497), .B1(n_1_674), .B2(n_1_603), .C1(n_1_656), 
      .C2(n_1_637), .ZN(n_1_496));
   INV_X1 i_1_688 (.A(n_1_498), .ZN(n_1_497));
   OAI22_X1 i_1_689 (.A1(n_1_664), .A2(n_1_628), .B1(n_1_652), .B2(n_1_600), 
      .ZN(n_1_498));
   OR3_X1 i_1_690 (.A1(n_1_718), .A2(n_1_499), .A3(n_1_514), .ZN(n_261));
   OR4_X1 i_1_691 (.A1(n_1_511), .A2(n_1_508), .A3(n_1_503), .A4(n_1_500), 
      .ZN(n_1_499));
   OAI221_X1 i_1_692 (.A(n_1_501), .B1(n_1_621), .B2(n_1_556), .C1(n_1_632), 
      .C2(n_1_541), .ZN(n_1_500));
   INV_X1 i_1_693 (.A(n_1_502), .ZN(n_1_501));
   OAI22_X1 i_1_694 (.A1(n_1_673), .A2(n_1_581), .B1(n_1_640), .B2(n_1_553), 
      .ZN(n_1_502));
   OAI221_X1 i_1_695 (.A(n_1_506), .B1(n_1_656), .B2(n_1_560), .C1(n_1_563), 
      .C2(n_1_504), .ZN(n_1_503));
   INV_X1 i_1_696 (.A(n_1_505), .ZN(n_1_504));
   NOR2_X1 i_1_697 (.A1(n_1_779), .A2(n_1_663), .ZN(n_1_505));
   INV_X1 i_1_698 (.A(n_1_507), .ZN(n_1_506));
   OAI22_X1 i_1_699 (.A1(n_1_603), .A2(n_1_531), .B1(n_1_612), .B2(n_1_566), 
      .ZN(n_1_507));
   OAI221_X1 i_1_700 (.A(n_1_509), .B1(n_1_599), .B2(n_1_550), .C1(n_1_652), 
      .C2(n_1_578), .ZN(n_1_508));
   INV_X1 i_1_701 (.A(n_1_510), .ZN(n_1_509));
   OAI22_X1 i_1_702 (.A1(n_1_608), .A2(n_1_538), .B1(n_1_681), .B2(n_1_584), 
      .ZN(n_1_510));
   OAI221_X1 i_1_703 (.A(n_1_512), .B1(n_1_687), .B2(n_1_547), .C1(n_1_617), 
      .C2(n_1_572), .ZN(n_1_511));
   INV_X1 i_1_704 (.A(n_1_513), .ZN(n_1_512));
   OAI22_X1 i_1_705 (.A1(n_1_667), .A2(n_1_575), .B1(n_1_628), .B2(n_1_534), 
      .ZN(n_1_513));
   OAI21_X1 i_1_706 (.A(n_1_689), .B1(n_1_728), .B2(n_1_515), .ZN(n_1_514));
   NOR3_X1 i_1_707 (.A1(n_1_662), .A2(n_1_517), .A3(n_1_644), .ZN(n_1_515));
   INV_X1 i_1_708 (.A(n_1_517), .ZN(n_1_516));
   NOR2_X1 i_1_709 (.A1(n_1_772), .A2(n_1_663), .ZN(n_1_517));
   OR4_X1 i_1_710 (.A1(n_1_521), .A2(n_1_518), .A3(n_1_524), .A4(n_1_585), 
      .ZN(n_262));
   OAI221_X1 i_1_711 (.A(n_1_519), .B1(n_1_678), .B2(n_1_603), .C1(n_1_687), 
      .C2(n_1_625), .ZN(n_1_518));
   INV_X1 i_1_712 (.A(n_1_520), .ZN(n_1_519));
   OAI22_X1 i_1_713 (.A1(n_1_681), .A2(n_1_674), .B1(n_1_664), .B2(n_1_652), 
      .ZN(n_1_520));
   OAI221_X1 i_1_714 (.A(n_1_522), .B1(n_1_684), .B2(n_1_632), .C1(n_1_656), 
      .C2(n_1_618), .ZN(n_1_521));
   INV_X1 i_1_715 (.A(n_1_523), .ZN(n_1_522));
   OAI22_X1 i_1_716 (.A1(n_1_673), .A2(n_1_629), .B1(n_1_640), .B2(n_1_605), 
      .ZN(n_1_523));
   OR4_X1 i_1_717 (.A1(n_1_528), .A2(n_1_527), .A3(n_1_526), .A4(n_1_525), 
      .ZN(n_1_524));
   OAI22_X1 i_1_718 (.A1(n_1_667), .A2(n_1_600), .B1(n_1_670), .B2(n_1_599), 
      .ZN(n_1_525));
   OAI21_X1 i_1_719 (.A(n_1_642), .B1(n_1_609), .B2(n_1_608), .ZN(n_1_526));
   OAI22_X1 i_1_720 (.A1(n_1_649), .A2(n_1_628), .B1(n_1_612), .B2(n_1_596), 
      .ZN(n_1_527));
   OAI22_X1 i_1_721 (.A1(n_1_653), .A2(n_1_617), .B1(n_1_637), .B2(n_1_621), 
      .ZN(n_1_528));
   OR3_X1 i_1_722 (.A1(n_1_569), .A2(n_1_529), .A3(n_1_585), .ZN(n_263));
   OR4_X1 i_1_723 (.A1(n_1_537), .A2(n_1_530), .A3(n_1_544), .A4(n_1_559), 
      .ZN(n_1_529));
   OAI22_X1 i_1_724 (.A1(n_1_652), .A2(n_1_534), .B1(n_1_681), .B2(n_1_531), 
      .ZN(n_1_530));
   INV_X1 i_1_725 (.A(n_1_532), .ZN(n_1_531));
   OAI221_X1 i_1_726 (.A(n_1_533), .B1(n_1_861), .B2(n_1_733), .C1(n_1_892), 
      .C2(n_1_734), .ZN(n_1_532));
   AOI22_X1 i_1_727 (.A1(a[1]), .A2(n_1_732), .B1(firstInputComplement[1]), 
      .B2(n_1_731), .ZN(n_1_533));
   INV_X1 i_1_728 (.A(n_1_535), .ZN(n_1_534));
   OAI221_X1 i_1_729 (.A(n_1_536), .B1(n_1_867), .B2(n_1_733), .C1(n_1_898), 
      .C2(n_1_734), .ZN(n_1_535));
   AOI22_X1 i_1_730 (.A1(a[7]), .A2(n_1_732), .B1(firstInputComplement[7]), 
      .B2(n_1_731), .ZN(n_1_536));
   OAI22_X1 i_1_731 (.A1(n_1_687), .A2(n_1_541), .B1(n_1_612), .B2(n_1_538), 
      .ZN(n_1_537));
   INV_X1 i_1_732 (.A(n_1_539), .ZN(n_1_538));
   OAI221_X1 i_1_733 (.A(n_1_540), .B1(n_1_879), .B2(n_1_733), .C1(n_1_910), 
      .C2(n_1_734), .ZN(n_1_539));
   AOI22_X1 i_1_734 (.A1(a[19]), .A2(n_1_732), .B1(firstInputComplement[19]), 
      .B2(n_1_731), .ZN(n_1_540));
   INV_X1 i_1_735 (.A(n_1_542), .ZN(n_1_541));
   OAI221_X1 i_1_736 (.A(n_1_543), .B1(n_1_871), .B2(n_1_733), .C1(n_1_902), 
      .C2(n_1_734), .ZN(n_1_542));
   AOI22_X1 i_1_737 (.A1(a[11]), .A2(n_1_732), .B1(firstInputComplement[11]), 
      .B2(n_1_731), .ZN(n_1_543));
   OAI221_X1 i_1_738 (.A(n_1_545), .B1(n_1_640), .B2(n_1_556), .C1(n_1_608), 
      .C2(n_1_553), .ZN(n_1_544));
   INV_X1 i_1_739 (.A(n_1_546), .ZN(n_1_545));
   OAI22_X1 i_1_740 (.A1(n_1_673), .A2(n_1_550), .B1(n_1_628), .B2(n_1_547), 
      .ZN(n_1_546));
   INV_X1 i_1_741 (.A(n_1_548), .ZN(n_1_547));
   OAI221_X1 i_1_742 (.A(n_1_549), .B1(n_1_869), .B2(n_1_733), .C1(n_1_900), 
      .C2(n_1_734), .ZN(n_1_548));
   AOI22_X1 i_1_743 (.A1(a[9]), .A2(n_1_732), .B1(firstInputComplement[9]), 
      .B2(n_1_731), .ZN(n_1_549));
   INV_X1 i_1_744 (.A(n_1_551), .ZN(n_1_550));
   OAI221_X1 i_1_745 (.A(n_1_552), .B1(n_1_875), .B2(n_1_733), .C1(n_1_906), 
      .C2(n_1_734), .ZN(n_1_551));
   AOI22_X1 i_1_746 (.A1(a[15]), .A2(n_1_732), .B1(firstInputComplement[15]), 
      .B2(n_1_731), .ZN(n_1_552));
   INV_X1 i_1_747 (.A(n_1_554), .ZN(n_1_553));
   OAI221_X1 i_1_748 (.A(n_1_555), .B1(n_1_881), .B2(n_1_733), .C1(n_1_912), 
      .C2(n_1_734), .ZN(n_1_554));
   AOI22_X1 i_1_749 (.A1(a[21]), .A2(n_1_732), .B1(firstInputComplement[21]), 
      .B2(n_1_731), .ZN(n_1_555));
   INV_X1 i_1_750 (.A(n_1_557), .ZN(n_1_556));
   OAI221_X1 i_1_751 (.A(n_1_558), .B1(n_1_883), .B2(n_1_733), .C1(n_1_914), 
      .C2(n_1_734), .ZN(n_1_557));
   AOI22_X1 i_1_752 (.A1(a[23]), .A2(n_1_732), .B1(firstInputComplement[23]), 
      .B2(n_1_731), .ZN(n_1_558));
   OAI222_X1 i_1_753 (.A1(n_1_617), .A2(n_1_563), .B1(n_1_621), .B2(n_1_560), 
      .C1(n_1_599), .C2(n_1_566), .ZN(n_1_559));
   INV_X1 i_1_754 (.A(n_1_561), .ZN(n_1_560));
   OAI221_X1 i_1_755 (.A(n_1_562), .B1(n_1_885), .B2(n_1_733), .C1(n_1_916), 
      .C2(n_1_734), .ZN(n_1_561));
   AOI22_X1 i_1_756 (.A1(a[25]), .A2(n_1_732), .B1(firstInputComplement[25]), 
      .B2(n_1_731), .ZN(n_1_562));
   INV_X1 i_1_757 (.A(n_1_564), .ZN(n_1_563));
   OAI221_X1 i_1_758 (.A(n_1_565), .B1(n_1_889), .B2(n_1_733), .C1(n_1_920), 
      .C2(n_1_734), .ZN(n_1_564));
   AOI22_X1 i_1_759 (.A1(a[29]), .A2(n_1_732), .B1(firstInputComplement[29]), 
      .B2(n_1_731), .ZN(n_1_565));
   INV_X1 i_1_760 (.A(n_1_567), .ZN(n_1_566));
   OAI221_X1 i_1_761 (.A(n_1_568), .B1(n_1_877), .B2(n_1_733), .C1(n_1_908), 
      .C2(n_1_734), .ZN(n_1_567));
   AOI22_X1 i_1_762 (.A1(a[17]), .A2(n_1_732), .B1(firstInputComplement[17]), 
      .B2(n_1_731), .ZN(n_1_568));
   OAI211_X1 i_1_763 (.A(n_1_642), .B(n_1_570), .C1(n_1_677), .C2(n_1_584), 
      .ZN(n_1_569));
   AOI221_X1 i_1_764 (.A(n_1_571), .B1(n_1_633), .B2(n_1_582), .C1(n_1_668), 
      .C2(n_1_579), .ZN(n_1_570));
   OAI22_X1 i_1_765 (.A1(n_1_603), .A2(n_1_575), .B1(n_1_656), .B2(n_1_572), 
      .ZN(n_1_571));
   INV_X1 i_1_766 (.A(n_1_573), .ZN(n_1_572));
   OAI221_X1 i_1_767 (.A(n_1_574), .B1(n_1_887), .B2(n_1_733), .C1(n_1_918), 
      .C2(n_1_734), .ZN(n_1_573));
   AOI22_X1 i_1_768 (.A1(a[27]), .A2(n_1_732), .B1(firstInputComplement[27]), 
      .B2(n_1_731), .ZN(n_1_574));
   INV_X1 i_1_769 (.A(n_1_576), .ZN(n_1_575));
   OAI221_X1 i_1_770 (.A(n_1_577), .B1(n_1_863), .B2(n_1_733), .C1(n_1_894), 
      .C2(n_1_734), .ZN(n_1_576));
   AOI22_X1 i_1_771 (.A1(a[3]), .A2(n_1_732), .B1(firstInputComplement[3]), 
      .B2(n_1_731), .ZN(n_1_577));
   INV_X1 i_1_772 (.A(n_1_579), .ZN(n_1_578));
   OAI221_X1 i_1_773 (.A(n_1_580), .B1(n_1_865), .B2(n_1_733), .C1(n_1_896), 
      .C2(n_1_734), .ZN(n_1_579));
   AOI22_X1 i_1_774 (.A1(a[5]), .A2(n_1_732), .B1(firstInputComplement[5]), 
      .B2(n_1_731), .ZN(n_1_580));
   INV_X1 i_1_775 (.A(n_1_582), .ZN(n_1_581));
   OAI221_X1 i_1_776 (.A(n_1_583), .B1(n_1_873), .B2(n_1_733), .C1(n_1_904), 
      .C2(n_1_734), .ZN(n_1_582));
   AOI22_X1 i_1_777 (.A1(a[13]), .A2(n_1_732), .B1(firstInputComplement[13]), 
      .B2(n_1_731), .ZN(n_1_583));
   OR2_X1 i_1_778 (.A1(n_1_859), .A2(n_1_744), .ZN(n_1_584));
   OR2_X1 i_1_779 (.A1(n_1_588), .A2(n_1_586), .ZN(n_1_585));
   OR2_X1 i_1_780 (.A1(n_1_938), .A2(n_1_587), .ZN(n_1_586));
   OR2_X1 i_1_781 (.A1(n_1_723), .A2(n_1_660), .ZN(n_1_587));
   OR2_X1 i_1_782 (.A1(n_1_591), .A2(n_1_589), .ZN(n_1_588));
   OR2_X1 i_1_783 (.A1(n_1_705), .A2(n_1_590), .ZN(n_1_589));
   NOR2_X1 i_1_784 (.A1(n_1_721), .A2(n_1_716), .ZN(n_1_590));
   OR2_X1 i_1_785 (.A1(n_1_691), .A2(n_1_592), .ZN(n_1_591));
   OAI21_X1 i_1_786 (.A(n_1_694), .B1(counter[2]), .B2(n_1_720), .ZN(n_1_592));
   NOR2_X1 i_1_787 (.A1(counter[2]), .A2(n_1_720), .ZN(n_1_593));
   OR3_X1 i_1_788 (.A1(n_1_658), .A2(n_1_594), .A3(n_1_688), .ZN(n_264));
   OR4_X1 i_1_789 (.A1(n_1_604), .A2(n_1_595), .A3(n_1_615), .A4(n_1_634), 
      .ZN(n_1_594));
   OAI22_X1 i_1_790 (.A1(n_1_603), .A2(n_1_600), .B1(n_1_599), .B2(n_1_596), 
      .ZN(n_1_595));
   INV_X1 i_1_791 (.A(n_1_597), .ZN(n_1_596));
   OAI221_X1 i_1_792 (.A(n_1_598), .B1(n_1_878), .B2(n_1_733), .C1(n_1_909), 
      .C2(n_1_734), .ZN(n_1_597));
   AOI22_X1 i_1_793 (.A1(a[18]), .A2(n_1_732), .B1(firstInputComplement[18]), 
      .B2(n_1_731), .ZN(n_1_598));
   OR2_X1 i_1_794 (.A1(n_1_714), .A2(n_1_613), .ZN(n_1_599));
   INV_X1 i_1_795 (.A(n_1_601), .ZN(n_1_600));
   OAI221_X1 i_1_796 (.A(n_1_602), .B1(n_1_864), .B2(n_1_733), .C1(n_1_895), 
      .C2(n_1_734), .ZN(n_1_601));
   AOI22_X1 i_1_797 (.A1(a[4]), .A2(n_1_732), .B1(firstInputComplement[4]), 
      .B2(n_1_731), .ZN(n_1_602));
   OR4_X1 i_1_798 (.A1(n_1_935), .A2(n_1_788), .A3(n_1_715), .A4(n_1_683), 
      .ZN(n_1_603));
   OAI22_X1 i_1_799 (.A1(n_1_612), .A2(n_1_609), .B1(n_1_608), .B2(n_1_605), 
      .ZN(n_1_604));
   INV_X1 i_1_800 (.A(n_1_606), .ZN(n_1_605));
   OAI221_X1 i_1_801 (.A(n_1_607), .B1(n_1_882), .B2(n_1_733), .C1(n_1_913), 
      .C2(n_1_734), .ZN(n_1_606));
   AOI22_X1 i_1_802 (.A1(a[22]), .A2(n_1_732), .B1(firstInputComplement[22]), 
      .B2(n_1_731), .ZN(n_1_607));
   OR3_X1 i_1_803 (.A1(n_1_937), .A2(n_1_786), .A3(n_1_614), .ZN(n_1_608));
   INV_X1 i_1_804 (.A(n_1_610), .ZN(n_1_609));
   OAI221_X1 i_1_805 (.A(n_1_611), .B1(n_1_880), .B2(n_1_733), .C1(n_1_911), 
      .C2(n_1_734), .ZN(n_1_610));
   AOI22_X1 i_1_806 (.A1(a[20]), .A2(n_1_732), .B1(firstInputComplement[20]), 
      .B2(n_1_731), .ZN(n_1_611));
   OR2_X1 i_1_807 (.A1(n_1_715), .A2(n_1_613), .ZN(n_1_612));
   NAND4_X1 i_1_808 (.A1(n_1_936), .A2(n_1_716), .A3(counter[4]), .A4(n_1_614), 
      .ZN(n_1_613));
   OAI21_X1 i_1_809 (.A(n_1_936), .B1(n_1_935), .B2(n_1_788), .ZN(n_1_614));
   OAI221_X1 i_1_810 (.A(n_1_623), .B1(n_1_621), .B2(n_1_618), .C1(n_1_728), 
      .C2(n_1_617), .ZN(n_1_615));
   INV_X1 i_1_811 (.A(n_1_617), .ZN(n_1_616));
   NAND3_X1 i_1_812 (.A1(counter[4]), .A2(n_1_786), .A3(n_1_788), .ZN(n_1_617));
   INV_X1 i_1_813 (.A(n_1_619), .ZN(n_1_618));
   OAI221_X1 i_1_814 (.A(n_1_620), .B1(n_1_886), .B2(n_1_733), .C1(n_1_917), 
      .C2(n_1_734), .ZN(n_1_619));
   AOI22_X1 i_1_815 (.A1(a[26]), .A2(n_1_732), .B1(firstInputComplement[26]), 
      .B2(n_1_731), .ZN(n_1_620));
   INV_X1 i_1_816 (.A(n_1_622), .ZN(n_1_621));
   NOR2_X1 i_1_817 (.A1(counter[0]), .A2(n_1_641), .ZN(n_1_622));
   INV_X1 i_1_818 (.A(n_1_624), .ZN(n_1_623));
   OAI22_X1 i_1_819 (.A1(n_1_632), .A2(n_1_629), .B1(n_1_628), .B2(n_1_625), 
      .ZN(n_1_624));
   INV_X1 i_1_820 (.A(n_1_626), .ZN(n_1_625));
   OAI221_X1 i_1_821 (.A(n_1_627), .B1(n_1_870), .B2(n_1_733), .C1(n_1_901), 
      .C2(n_1_734), .ZN(n_1_626));
   AOI22_X1 i_1_822 (.A1(a[10]), .A2(n_1_732), .B1(firstInputComplement[10]), 
      .B2(n_1_731), .ZN(n_1_627));
   OR2_X1 i_1_823 (.A1(n_1_727), .A2(n_1_683), .ZN(n_1_628));
   INV_X1 i_1_824 (.A(n_1_630), .ZN(n_1_629));
   OAI221_X1 i_1_825 (.A(n_1_631), .B1(n_1_874), .B2(n_1_733), .C1(n_1_905), 
      .C2(n_1_734), .ZN(n_1_630));
   AOI22_X1 i_1_826 (.A1(a[14]), .A2(n_1_732), .B1(firstInputComplement[14]), 
      .B2(n_1_731), .ZN(n_1_631));
   INV_X1 i_1_827 (.A(n_1_633), .ZN(n_1_632));
   NOR3_X1 i_1_828 (.A1(counter[2]), .A2(n_1_787), .A3(n_1_683), .ZN(n_1_633));
   OAI221_X1 i_1_829 (.A(n_1_635), .B1(n_1_656), .B2(n_1_653), .C1(n_1_652), 
      .C2(n_1_649), .ZN(n_1_634));
   INV_X1 i_1_830 (.A(n_1_636), .ZN(n_1_635));
   OAI21_X1 i_1_831 (.A(n_1_642), .B1(n_1_640), .B2(n_1_637), .ZN(n_1_636));
   INV_X1 i_1_832 (.A(n_1_638), .ZN(n_1_637));
   OAI221_X1 i_1_833 (.A(n_1_639), .B1(n_1_884), .B2(n_1_733), .C1(n_1_915), 
      .C2(n_1_734), .ZN(n_1_638));
   AOI22_X1 i_1_834 (.A1(a[24]), .A2(n_1_732), .B1(firstInputComplement[24]), 
      .B2(n_1_731), .ZN(n_1_639));
   OR2_X1 i_1_835 (.A1(n_1_933), .A2(n_1_641), .ZN(n_1_640));
   NAND3_X1 i_1_836 (.A1(counter[4]), .A2(n_1_786), .A3(counter[1]), .ZN(n_1_641));
   OAI21_X1 i_1_837 (.A(n_1_729), .B1(n_1_644), .B2(n_1_643), .ZN(n_1_642));
   NOR3_X1 i_1_838 (.A1(counter[4]), .A2(n_1_714), .A3(n_1_936), .ZN(n_1_643));
   NAND2_X1 i_1_839 (.A1(n_1_647), .A2(n_1_645), .ZN(n_1_644));
   INV_X1 i_1_840 (.A(n_1_646), .ZN(n_1_645));
   NOR3_X1 i_1_841 (.A1(n_1_935), .A2(n_1_787), .A3(n_1_726), .ZN(n_1_646));
   INV_X1 i_1_842 (.A(n_1_648), .ZN(n_1_647));
   NOR3_X1 i_1_843 (.A1(counter[4]), .A2(n_1_774), .A3(n_1_779), .ZN(n_1_648));
   INV_X1 i_1_844 (.A(n_1_650), .ZN(n_1_649));
   OAI221_X1 i_1_845 (.A(n_1_651), .B1(n_1_868), .B2(n_1_733), .C1(n_1_899), 
      .C2(n_1_734), .ZN(n_1_650));
   AOI22_X1 i_1_846 (.A1(a[8]), .A2(n_1_732), .B1(firstInputComplement[8]), 
      .B2(n_1_731), .ZN(n_1_651));
   OR3_X1 i_1_847 (.A1(counter[2]), .A2(n_1_717), .A3(n_1_683), .ZN(n_1_652));
   INV_X1 i_1_848 (.A(n_1_654), .ZN(n_1_653));
   OAI221_X1 i_1_849 (.A(n_1_655), .B1(n_1_888), .B2(n_1_733), .C1(n_1_919), 
      .C2(n_1_734), .ZN(n_1_654));
   AOI22_X1 i_1_850 (.A1(a[28]), .A2(n_1_732), .B1(firstInputComplement[28]), 
      .B2(n_1_731), .ZN(n_1_655));
   NAND2_X1 i_1_851 (.A1(counter[0]), .A2(n_1_657), .ZN(n_1_656));
   NOR4_X1 i_1_852 (.A1(counter[3]), .A2(counter[2]), .A3(n_1_937), .A4(
      counter[1]), .ZN(n_1_657));
   OAI221_X1 i_1_853 (.A(n_1_659), .B1(n_1_687), .B2(n_1_684), .C1(n_1_681), 
      .C2(n_1_678), .ZN(n_1_658));
   AOI211_X1 i_1_854 (.A(n_1_660), .B(n_1_669), .C1(n_1_668), .C2(n_1_665), 
      .ZN(n_1_659));
   NOR2_X1 i_1_855 (.A1(n_1_728), .A2(n_1_661), .ZN(n_1_660));
   INV_X1 i_1_856 (.A(n_1_662), .ZN(n_1_661));
   NOR2_X1 i_1_857 (.A1(n_1_763), .A2(n_1_663), .ZN(n_1_662));
   NAND2_X1 i_1_858 (.A1(n_1_937), .A2(n_1_778), .ZN(n_1_663));
   INV_X1 i_1_859 (.A(n_1_665), .ZN(n_1_664));
   OAI221_X1 i_1_860 (.A(n_1_666), .B1(n_1_866), .B2(n_1_733), .C1(n_1_897), 
      .C2(n_1_734), .ZN(n_1_665));
   AOI22_X1 i_1_861 (.A1(a[6]), .A2(n_1_732), .B1(firstInputComplement[6]), 
      .B2(n_1_731), .ZN(n_1_666));
   INV_X1 i_1_862 (.A(n_1_668), .ZN(n_1_667));
   NOR3_X1 i_1_863 (.A1(n_1_935), .A2(n_1_787), .A3(n_1_683), .ZN(n_1_668));
   OAI22_X1 i_1_864 (.A1(n_1_677), .A2(n_1_674), .B1(n_1_673), .B2(n_1_670), 
      .ZN(n_1_669));
   INV_X1 i_1_865 (.A(n_1_671), .ZN(n_1_670));
   OAI221_X1 i_1_866 (.A(n_1_672), .B1(n_1_876), .B2(n_1_733), .C1(n_1_907), 
      .C2(n_1_734), .ZN(n_1_671));
   AOI22_X1 i_1_867 (.A1(a[16]), .A2(n_1_732), .B1(firstInputComplement[16]), 
      .B2(n_1_731), .ZN(n_1_672));
   NAND3_X1 i_1_868 (.A1(counter[4]), .A2(n_1_780), .A3(n_1_777), .ZN(n_1_673));
   INV_X1 i_1_869 (.A(n_1_675), .ZN(n_1_674));
   OAI221_X1 i_1_870 (.A(n_1_676), .B1(n_1_891), .B2(n_1_734), .C1(n_1_860), 
      .C2(n_1_733), .ZN(n_1_675));
   OAI21_X1 i_1_871 (.A(a[0]), .B1(n_1_732), .B2(n_1_731), .ZN(n_1_676));
   NAND2_X1 i_1_872 (.A1(counter[0]), .A2(n_1_682), .ZN(n_1_677));
   INV_X1 i_1_873 (.A(n_1_679), .ZN(n_1_678));
   OAI221_X1 i_1_874 (.A(n_1_680), .B1(n_1_862), .B2(n_1_733), .C1(n_1_893), 
      .C2(n_1_734), .ZN(n_1_679));
   AOI22_X1 i_1_875 (.A1(a[2]), .A2(n_1_732), .B1(firstInputComplement[2]), 
      .B2(n_1_731), .ZN(n_1_680));
   NAND2_X1 i_1_876 (.A1(n_1_717), .A2(n_1_682), .ZN(n_1_681));
   NOR2_X1 i_1_877 (.A1(n_1_714), .A2(n_1_683), .ZN(n_1_682));
   NAND2_X1 i_1_878 (.A1(counter[4]), .A2(counter[3]), .ZN(n_1_683));
   INV_X1 i_1_879 (.A(n_1_685), .ZN(n_1_684));
   OAI221_X1 i_1_880 (.A(n_1_686), .B1(n_1_872), .B2(n_1_733), .C1(n_1_903), 
      .C2(n_1_734), .ZN(n_1_685));
   AOI22_X1 i_1_881 (.A1(a[12]), .A2(n_1_732), .B1(firstInputComplement[12]), 
      .B2(n_1_731), .ZN(n_1_686));
   OR4_X1 i_1_882 (.A1(n_1_774), .A2(n_1_763), .A3(n_1_937), .A4(n_1_786), 
      .ZN(n_1_687));
   OR3_X1 i_1_883 (.A1(n_1_700), .A2(n_1_690), .A3(n_1_718), .ZN(n_1_688));
   NOR2_X1 i_1_884 (.A1(n_1_700), .A2(n_1_690), .ZN(n_1_689));
   OAI21_X1 i_1_885 (.A(n_1_694), .B1(n_1_728), .B2(n_1_692), .ZN(n_1_690));
   NOR2_X1 i_1_886 (.A1(n_1_728), .A2(n_1_692), .ZN(n_1_691));
   OR2_X1 i_1_887 (.A1(n_1_772), .A2(n_1_709), .ZN(n_1_692));
   INV_X1 i_1_888 (.A(n_1_694), .ZN(n_1_693));
   NOR2_X1 i_1_889 (.A1(n_1_699), .A2(n_1_695), .ZN(n_1_694));
   NOR2_X1 i_1_890 (.A1(n_1_728), .A2(n_1_696), .ZN(n_1_695));
   INV_X1 i_1_891 (.A(n_1_697), .ZN(n_1_696));
   NOR2_X1 i_1_892 (.A1(n_1_763), .A2(n_1_709), .ZN(n_1_697));
   INV_X1 i_1_893 (.A(n_1_699), .ZN(n_1_698));
   NOR2_X1 i_1_894 (.A1(n_1_785), .A2(n_1_728), .ZN(n_1_699));
   OR2_X1 i_1_895 (.A1(n_1_705), .A2(n_1_938), .ZN(n_1_700));
   INV_X1 i_1_896 (.A(n_1_702), .ZN(n_1_701));
   NOR3_X1 i_1_897 (.A1(n_1_774), .A2(n_1_763), .A3(counter[4]), .ZN(n_1_702));
   NOR2_X1 i_1_898 (.A1(n_1_728), .A2(n_1_704), .ZN(n_1_703));
   NAND4_X1 i_1_899 (.A1(n_1_937), .A2(counter[3]), .A3(n_1_935), .A4(n_1_788), 
      .ZN(n_1_704));
   OAI21_X1 i_1_900 (.A(n_1_710), .B1(n_1_728), .B2(n_1_707), .ZN(n_1_705));
   NOR2_X1 i_1_901 (.A1(n_1_728), .A2(n_1_707), .ZN(n_1_706));
   INV_X1 i_1_902 (.A(n_1_708), .ZN(n_1_707));
   NOR2_X1 i_1_903 (.A1(n_1_779), .A2(n_1_709), .ZN(n_1_708));
   NAND3_X1 i_1_904 (.A1(n_1_937), .A2(n_1_936), .A3(n_1_934), .ZN(n_1_709));
   INV_X1 i_1_905 (.A(n_1_711), .ZN(n_1_710));
   NOR2_X1 i_1_906 (.A1(n_1_728), .A2(n_1_713), .ZN(n_1_711));
   INV_X1 i_1_907 (.A(n_1_713), .ZN(n_1_712));
   NAND4_X1 i_1_908 (.A1(n_1_936), .A2(n_1_716), .A3(n_1_937), .A4(n_1_715), 
      .ZN(n_1_713));
   INV_X1 i_1_909 (.A(n_1_715), .ZN(n_1_714));
   NOR2_X1 i_1_910 (.A1(n_1_935), .A2(n_1_934), .ZN(n_1_715));
   NAND3_X1 i_1_911 (.A1(counter[1]), .A2(counter[0]), .A3(counter[2]), .ZN(
      n_1_716));
   NAND2_X1 i_1_912 (.A1(counter[1]), .A2(counter[0]), .ZN(n_1_717));
   OR2_X1 i_1_913 (.A1(n_1_723), .A2(n_1_719), .ZN(n_1_718));
   NOR2_X1 i_1_914 (.A1(n_1_773), .A2(n_1_720), .ZN(n_1_719));
   OR2_X1 i_1_915 (.A1(n_1_934), .A2(n_1_721), .ZN(n_1_720));
   NAND3_X1 i_1_916 (.A1(n_1_937), .A2(n_1_936), .A3(n_1_729), .ZN(n_1_721));
   NAND2_X1 i_1_917 (.A1(n_1_937), .A2(n_1_936), .ZN(n_1_722));
   NOR2_X1 i_1_918 (.A1(n_1_728), .A2(n_1_724), .ZN(n_1_723));
   INV_X1 i_1_919 (.A(n_1_725), .ZN(n_1_724));
   NOR2_X1 i_1_920 (.A1(n_1_727), .A2(n_1_726), .ZN(n_1_725));
   NAND2_X1 i_1_921 (.A1(n_1_937), .A2(counter[3]), .ZN(n_1_726));
   NAND3_X1 i_1_922 (.A1(n_1_935), .A2(n_1_933), .A3(counter[1]), .ZN(n_1_727));
   INV_X1 i_1_923 (.A(n_1_729), .ZN(n_1_728));
   OAI221_X1 i_1_924 (.A(n_1_730), .B1(n_1_890), .B2(n_1_733), .C1(n_1_921), 
      .C2(n_1_734), .ZN(n_1_729));
   AOI22_X1 i_1_925 (.A1(a[30]), .A2(n_1_732), .B1(firstInputComplement[30]), 
      .B2(n_1_731), .ZN(n_1_730));
   NOR2_X1 i_1_926 (.A1(n_1_745), .A2(n_1_736), .ZN(n_1_731));
   NOR2_X1 i_1_927 (.A1(n_1_746), .A2(n_1_735), .ZN(n_1_732));
   OR2_X1 i_1_928 (.A1(n_1_744), .A2(n_1_735), .ZN(n_1_733));
   OR2_X1 i_1_929 (.A1(n_1_744), .A2(n_1_736), .ZN(n_1_734));
   INV_X1 i_1_930 (.A(n_1_736), .ZN(n_1_735));
   NOR3_X1 i_1_931 (.A1(n_1_741), .A2(n_1_738), .A3(n_1_737), .ZN(n_1_736));
   OAI22_X1 i_1_932 (.A1(n_1_760), .A2(n_1_750), .B1(n_1_772), .B2(n_1_754), 
      .ZN(n_1_737));
   OAI22_X1 i_1_933 (.A1(n_1_774), .A2(n_1_740), .B1(n_1_768), .B2(n_1_739), 
      .ZN(n_1_738));
   AOI22_X1 i_1_934 (.A1(b[11]), .A2(n_1_780), .B1(b[3]), .B2(n_1_764), .ZN(
      n_1_739));
   AOI22_X1 i_1_935 (.A1(b[19]), .A2(n_1_764), .B1(b[27]), .B2(n_1_780), 
      .ZN(n_1_740));
   OAI22_X1 i_1_936 (.A1(n_1_763), .A2(n_1_743), .B1(n_1_779), .B2(n_1_742), 
      .ZN(n_1_741));
   AOI22_X1 i_1_937 (.A1(b[15]), .A2(n_1_777), .B1(b[31]), .B2(n_1_778), 
      .ZN(n_1_742));
   AOI22_X1 i_1_938 (.A1(b[23]), .A2(n_1_778), .B1(b[7]), .B2(n_1_777), .ZN(
      n_1_743));
   NAND2_X1 i_1_939 (.A1(n_1_746), .A2(n_1_745), .ZN(n_1_744));
   OR2_X1 i_1_940 (.A1(n_1_757), .A2(n_1_747), .ZN(n_1_745));
   NAND2_X1 i_1_941 (.A1(n_1_757), .A2(n_1_747), .ZN(n_1_746));
   OAI221_X1 i_1_942 (.A(n_1_752), .B1(n_1_763), .B2(n_1_750), .C1(n_1_772), 
      .C2(n_1_748), .ZN(n_1_747));
   AOI221_X1 i_1_943 (.A(n_1_749), .B1(b[11]), .B2(n_1_777), .C1(b[27]), 
      .C2(n_1_778), .ZN(n_1_748));
   OAI22_X1 i_1_944 (.A1(n_1_931), .A2(n_1_774), .B1(n_1_926), .B2(n_1_768), 
      .ZN(n_1_749));
   AOI221_X1 i_1_945 (.A(n_1_751), .B1(b[5]), .B2(n_1_777), .C1(b[21]), .C2(
      n_1_778), .ZN(n_1_750));
   OAI22_X1 i_1_946 (.A1(n_1_924), .A2(n_1_768), .B1(n_1_929), .B2(n_1_774), 
      .ZN(n_1_751));
   INV_X1 i_1_947 (.A(n_1_753), .ZN(n_1_752));
   OAI22_X1 i_1_948 (.A1(n_1_760), .A2(n_1_756), .B1(n_1_779), .B2(n_1_754), 
      .ZN(n_1_753));
   AOI221_X1 i_1_949 (.A(n_1_755), .B1(b[29]), .B2(n_1_778), .C1(b[13]), 
      .C2(n_1_777), .ZN(n_1_754));
   OAI22_X1 i_1_950 (.A1(n_1_927), .A2(n_1_768), .B1(n_1_932), .B2(n_1_774), 
      .ZN(n_1_755));
   AOI222_X1 i_1_951 (.A1(b[3]), .A2(n_1_777), .B1(b[15]), .B2(n_1_775), 
      .C1(b[19]), .C2(n_1_778), .ZN(n_1_756));
   OAI221_X1 i_1_952 (.A(n_1_765), .B1(n_1_763), .B2(n_1_761), .C1(n_1_760), 
      .C2(n_1_758), .ZN(n_1_757));
   AOI221_X1 i_1_953 (.A(n_1_759), .B1(b[20]), .B2(n_1_778), .C1(b[4]), .C2(
      n_1_777), .ZN(n_1_758));
   OAI22_X1 i_1_954 (.A1(n_1_923), .A2(n_1_768), .B1(n_1_928), .B2(n_1_774), 
      .ZN(n_1_759));
   NAND2_X1 i_1_955 (.A1(n_1_935), .A2(n_1_933), .ZN(n_1_760));
   AOI221_X1 i_1_956 (.A(n_1_762), .B1(b[6]), .B2(n_1_777), .C1(b[22]), .C2(
      n_1_778), .ZN(n_1_761));
   OAI22_X1 i_1_957 (.A1(n_1_930), .A2(n_1_774), .B1(n_1_925), .B2(n_1_768), 
      .ZN(n_1_762));
   INV_X1 i_1_958 (.A(n_1_764), .ZN(n_1_763));
   NOR2_X1 i_1_959 (.A1(counter[2]), .A2(n_1_933), .ZN(n_1_764));
   NOR2_X1 i_1_960 (.A1(n_1_770), .A2(n_1_766), .ZN(n_1_765));
   OAI22_X1 i_1_961 (.A1(n_1_772), .A2(n_1_769), .B1(n_1_768), .B2(n_1_767), 
      .ZN(n_1_766));
   AOI22_X1 i_1_962 (.A1(b[10]), .A2(n_1_780), .B1(b[8]), .B2(n_1_773), .ZN(
      n_1_767));
   NAND2_X1 i_1_963 (.A1(n_1_936), .A2(n_1_934), .ZN(n_1_768));
   AOI22_X1 i_1_964 (.A1(b[12]), .A2(n_1_777), .B1(b[28]), .B2(n_1_778), 
      .ZN(n_1_769));
   OAI22_X1 i_1_965 (.A1(n_1_779), .A2(n_1_776), .B1(n_1_774), .B2(n_1_771), 
      .ZN(n_1_770));
   AOI22_X1 i_1_966 (.A1(b[24]), .A2(n_1_773), .B1(b[26]), .B2(n_1_780), 
      .ZN(n_1_771));
   INV_X1 i_1_967 (.A(n_1_773), .ZN(n_1_772));
   NOR2_X1 i_1_968 (.A1(n_1_935), .A2(counter[0]), .ZN(n_1_773));
   INV_X1 i_1_969 (.A(n_1_775), .ZN(n_1_774));
   NOR2_X1 i_1_970 (.A1(n_1_936), .A2(counter[1]), .ZN(n_1_775));
   AOI22_X1 i_1_971 (.A1(b[30]), .A2(n_1_778), .B1(b[14]), .B2(n_1_777), 
      .ZN(n_1_776));
   NOR2_X1 i_1_972 (.A1(counter[3]), .A2(n_1_934), .ZN(n_1_777));
   NOR2_X1 i_1_973 (.A1(n_1_936), .A2(n_1_934), .ZN(n_1_778));
   INV_X1 i_1_974 (.A(n_1_780), .ZN(n_1_779));
   NOR2_X1 i_1_975 (.A1(n_1_935), .A2(n_1_933), .ZN(n_1_780));
   NOR3_X1 i_1_976 (.A1(n_1_922), .A2(reset), .A3(resetReg), .ZN(n_265));
   OAI21_X1 i_1_977 (.A(n_1_782), .B1(n_1_789), .B2(n_1_781), .ZN(n_266));
   NOR2_X1 i_1_978 (.A1(n_1_922), .A2(n_1_785), .ZN(n_1_781));
   INV_X1 i_1_979 (.A(n_1_782), .ZN(n_267));
   OAI21_X1 i_1_980 (.A(en), .B1(reset), .B2(resetReg), .ZN(n_1_782));
   OAI21_X1 i_1_981 (.A(en), .B1(n_1_789), .B2(n_1_783), .ZN(n_268));
   OR3_X1 i_1_982 (.A1(reset), .A2(resetReg), .A3(n_1_784), .ZN(n_1_783));
   INV_X1 i_1_983 (.A(n_1_785), .ZN(n_1_784));
   NAND3_X1 i_1_984 (.A1(n_1_788), .A2(n_1_786), .A3(n_1_937), .ZN(n_1_785));
   NOR2_X1 i_1_985 (.A1(counter[3]), .A2(counter[2]), .ZN(n_1_786));
   INV_X1 i_1_986 (.A(n_1_788), .ZN(n_1_787));
   NOR2_X1 i_1_987 (.A1(counter[1]), .A2(counter[0]), .ZN(n_1_788));
   OR2_X1 i_1_988 (.A1(n_1_791), .A2(n_1_790), .ZN(n_1_789));
   NAND4_X1 i_1_989 (.A1(counter[0]), .A2(n_1_794), .A3(n_1_793), .A4(n_1_792), 
      .ZN(n_1_790));
   XOR2_X1 i_1_990 (.A(n_1_937), .B(n_1_2), .Z(n_1_791));
   INV_X1 i_1_991 (.A(n_1_5), .ZN(n_1_792));
   INV_X1 i_1_992 (.A(n_1_4), .ZN(n_1_793));
   INV_X1 i_1_993 (.A(n_1_3), .ZN(n_1_794));
   INV_X1 i_1_994 (.A(n_3), .ZN(n_1_795));
   INV_X1 i_1_995 (.A(n_4), .ZN(n_1_796));
   INV_X1 i_1_996 (.A(n_5), .ZN(n_1_797));
   INV_X1 i_1_997 (.A(n_6), .ZN(n_1_798));
   INV_X1 i_1_998 (.A(n_7), .ZN(n_1_799));
   INV_X1 i_1_999 (.A(n_8), .ZN(n_1_800));
   INV_X1 i_1_1000 (.A(n_9), .ZN(n_1_801));
   INV_X1 i_1_1001 (.A(n_10), .ZN(n_1_802));
   INV_X1 i_1_1002 (.A(n_11), .ZN(n_1_803));
   INV_X1 i_1_1003 (.A(n_12), .ZN(n_1_804));
   INV_X1 i_1_1004 (.A(n_13), .ZN(n_1_805));
   INV_X1 i_1_1005 (.A(n_14), .ZN(n_1_806));
   INV_X1 i_1_1006 (.A(n_15), .ZN(n_1_807));
   INV_X1 i_1_1007 (.A(n_16), .ZN(n_1_808));
   INV_X1 i_1_1008 (.A(n_17), .ZN(n_1_809));
   INV_X1 i_1_1009 (.A(n_18), .ZN(n_1_810));
   INV_X1 i_1_1010 (.A(n_19), .ZN(n_1_811));
   INV_X1 i_1_1011 (.A(n_20), .ZN(n_1_812));
   INV_X1 i_1_1012 (.A(n_21), .ZN(n_1_813));
   INV_X1 i_1_1013 (.A(n_22), .ZN(n_1_814));
   INV_X1 i_1_1014 (.A(n_23), .ZN(n_1_815));
   INV_X1 i_1_1015 (.A(n_24), .ZN(n_1_816));
   INV_X1 i_1_1016 (.A(n_25), .ZN(n_1_817));
   INV_X1 i_1_1017 (.A(n_26), .ZN(n_1_818));
   INV_X1 i_1_1018 (.A(n_27), .ZN(n_1_819));
   INV_X1 i_1_1019 (.A(n_28), .ZN(n_1_820));
   INV_X1 i_1_1020 (.A(n_29), .ZN(n_1_821));
   INV_X1 i_1_1021 (.A(n_30), .ZN(n_1_822));
   INV_X1 i_1_1022 (.A(n_31), .ZN(n_1_823));
   INV_X1 i_1_1023 (.A(n_32), .ZN(n_1_824));
   INV_X1 i_1_1024 (.A(n_33), .ZN(n_1_825));
   INV_X1 i_1_1025 (.A(n_34), .ZN(n_1_826));
   INV_X1 i_1_1026 (.A(n_35), .ZN(n_1_827));
   INV_X1 i_1_1027 (.A(n_36), .ZN(n_1_828));
   INV_X1 i_1_1028 (.A(n_37), .ZN(n_1_829));
   INV_X1 i_1_1029 (.A(n_38), .ZN(n_1_830));
   INV_X1 i_1_1030 (.A(n_39), .ZN(n_1_831));
   INV_X1 i_1_1031 (.A(n_40), .ZN(n_1_832));
   INV_X1 i_1_1032 (.A(n_41), .ZN(n_1_833));
   INV_X1 i_1_1033 (.A(n_42), .ZN(n_1_834));
   INV_X1 i_1_1034 (.A(n_43), .ZN(n_1_835));
   INV_X1 i_1_1035 (.A(n_44), .ZN(n_1_836));
   INV_X1 i_1_1036 (.A(n_45), .ZN(n_1_837));
   INV_X1 i_1_1037 (.A(n_46), .ZN(n_1_838));
   INV_X1 i_1_1038 (.A(n_47), .ZN(n_1_839));
   INV_X1 i_1_1039 (.A(n_48), .ZN(n_1_840));
   INV_X1 i_1_1040 (.A(n_49), .ZN(n_1_841));
   INV_X1 i_1_1041 (.A(n_50), .ZN(n_1_842));
   INV_X1 i_1_1042 (.A(n_51), .ZN(n_1_843));
   INV_X1 i_1_1043 (.A(n_52), .ZN(n_1_844));
   INV_X1 i_1_1044 (.A(n_53), .ZN(n_1_845));
   INV_X1 i_1_1045 (.A(n_54), .ZN(n_1_846));
   INV_X1 i_1_1046 (.A(n_55), .ZN(n_1_847));
   INV_X1 i_1_1047 (.A(n_56), .ZN(n_1_848));
   INV_X1 i_1_1048 (.A(n_57), .ZN(n_1_849));
   INV_X1 i_1_1049 (.A(n_58), .ZN(n_1_850));
   INV_X1 i_1_1050 (.A(n_59), .ZN(n_1_851));
   INV_X1 i_1_1051 (.A(n_60), .ZN(n_1_852));
   INV_X1 i_1_1052 (.A(n_61), .ZN(n_1_853));
   INV_X1 i_1_1053 (.A(n_62), .ZN(n_1_854));
   INV_X1 i_1_1054 (.A(n_63), .ZN(n_1_855));
   INV_X1 i_1_1055 (.A(n_64), .ZN(n_1_856));
   INV_X1 i_1_1056 (.A(n_65), .ZN(n_1_857));
   INV_X1 i_1_1057 (.A(n_66), .ZN(n_1_858));
   INV_X1 i_1_1058 (.A(a[0]), .ZN(n_1_859));
   INV_X1 i_1_1059 (.A(a[1]), .ZN(n_1_860));
   INV_X1 i_1_1060 (.A(a[2]), .ZN(n_1_861));
   INV_X1 i_1_1061 (.A(a[3]), .ZN(n_1_862));
   INV_X1 i_1_1062 (.A(a[4]), .ZN(n_1_863));
   INV_X1 i_1_1063 (.A(a[5]), .ZN(n_1_864));
   INV_X1 i_1_1064 (.A(a[6]), .ZN(n_1_865));
   INV_X1 i_1_1065 (.A(a[7]), .ZN(n_1_866));
   INV_X1 i_1_1066 (.A(a[8]), .ZN(n_1_867));
   INV_X1 i_1_1067 (.A(a[9]), .ZN(n_1_868));
   INV_X1 i_1_1068 (.A(a[10]), .ZN(n_1_869));
   INV_X1 i_1_1069 (.A(a[11]), .ZN(n_1_870));
   INV_X1 i_1_1070 (.A(a[12]), .ZN(n_1_871));
   INV_X1 i_1_1071 (.A(a[13]), .ZN(n_1_872));
   INV_X1 i_1_1072 (.A(a[14]), .ZN(n_1_873));
   INV_X1 i_1_1073 (.A(a[15]), .ZN(n_1_874));
   INV_X1 i_1_1074 (.A(a[16]), .ZN(n_1_875));
   INV_X1 i_1_1075 (.A(a[17]), .ZN(n_1_876));
   INV_X1 i_1_1076 (.A(a[18]), .ZN(n_1_877));
   INV_X1 i_1_1077 (.A(a[19]), .ZN(n_1_878));
   INV_X1 i_1_1078 (.A(a[20]), .ZN(n_1_879));
   INV_X1 i_1_1079 (.A(a[21]), .ZN(n_1_880));
   INV_X1 i_1_1080 (.A(a[22]), .ZN(n_1_881));
   INV_X1 i_1_1081 (.A(a[23]), .ZN(n_1_882));
   INV_X1 i_1_1082 (.A(a[24]), .ZN(n_1_883));
   INV_X1 i_1_1083 (.A(a[25]), .ZN(n_1_884));
   INV_X1 i_1_1084 (.A(a[26]), .ZN(n_1_885));
   INV_X1 i_1_1085 (.A(a[27]), .ZN(n_1_886));
   INV_X1 i_1_1086 (.A(a[28]), .ZN(n_1_887));
   INV_X1 i_1_1087 (.A(a[29]), .ZN(n_1_888));
   INV_X1 i_1_1088 (.A(a[30]), .ZN(n_1_889));
   INV_X1 i_1_1089 (.A(a[31]), .ZN(n_1_890));
   INV_X1 i_1_1090 (.A(firstInputComplement[1]), .ZN(n_1_891));
   INV_X1 i_1_1091 (.A(firstInputComplement[2]), .ZN(n_1_892));
   INV_X1 i_1_1092 (.A(firstInputComplement[3]), .ZN(n_1_893));
   INV_X1 i_1_1093 (.A(firstInputComplement[4]), .ZN(n_1_894));
   INV_X1 i_1_1094 (.A(firstInputComplement[5]), .ZN(n_1_895));
   INV_X1 i_1_1095 (.A(firstInputComplement[6]), .ZN(n_1_896));
   INV_X1 i_1_1096 (.A(firstInputComplement[7]), .ZN(n_1_897));
   INV_X1 i_1_1097 (.A(firstInputComplement[8]), .ZN(n_1_898));
   INV_X1 i_1_1098 (.A(firstInputComplement[9]), .ZN(n_1_899));
   INV_X1 i_1_1099 (.A(firstInputComplement[10]), .ZN(n_1_900));
   INV_X1 i_1_1100 (.A(firstInputComplement[11]), .ZN(n_1_901));
   INV_X1 i_1_1101 (.A(firstInputComplement[12]), .ZN(n_1_902));
   INV_X1 i_1_1102 (.A(firstInputComplement[13]), .ZN(n_1_903));
   INV_X1 i_1_1103 (.A(firstInputComplement[14]), .ZN(n_1_904));
   INV_X1 i_1_1104 (.A(firstInputComplement[15]), .ZN(n_1_905));
   INV_X1 i_1_1105 (.A(firstInputComplement[16]), .ZN(n_1_906));
   INV_X1 i_1_1106 (.A(firstInputComplement[17]), .ZN(n_1_907));
   INV_X1 i_1_1107 (.A(firstInputComplement[18]), .ZN(n_1_908));
   INV_X1 i_1_1108 (.A(firstInputComplement[19]), .ZN(n_1_909));
   INV_X1 i_1_1109 (.A(firstInputComplement[20]), .ZN(n_1_910));
   INV_X1 i_1_1110 (.A(firstInputComplement[21]), .ZN(n_1_911));
   INV_X1 i_1_1111 (.A(firstInputComplement[22]), .ZN(n_1_912));
   INV_X1 i_1_1112 (.A(firstInputComplement[23]), .ZN(n_1_913));
   INV_X1 i_1_1113 (.A(firstInputComplement[24]), .ZN(n_1_914));
   INV_X1 i_1_1114 (.A(firstInputComplement[25]), .ZN(n_1_915));
   INV_X1 i_1_1115 (.A(firstInputComplement[26]), .ZN(n_1_916));
   INV_X1 i_1_1116 (.A(firstInputComplement[27]), .ZN(n_1_917));
   INV_X1 i_1_1117 (.A(firstInputComplement[28]), .ZN(n_1_918));
   INV_X1 i_1_1118 (.A(firstInputComplement[29]), .ZN(n_1_919));
   INV_X1 i_1_1119 (.A(firstInputComplement[30]), .ZN(n_1_920));
   INV_X1 i_1_1120 (.A(firstInputComplement[31]), .ZN(n_1_921));
   INV_X1 i_1_1121 (.A(en), .ZN(n_1_922));
   INV_X1 i_1_1122 (.A(b[0]), .ZN(n_1_923));
   INV_X1 i_1_1123 (.A(b[1]), .ZN(n_1_924));
   INV_X1 i_1_1124 (.A(b[2]), .ZN(n_1_925));
   INV_X1 i_1_1125 (.A(b[7]), .ZN(n_1_926));
   INV_X1 i_1_1126 (.A(b[9]), .ZN(n_1_927));
   INV_X1 i_1_1127 (.A(b[16]), .ZN(n_1_928));
   INV_X1 i_1_1128 (.A(b[17]), .ZN(n_1_929));
   INV_X1 i_1_1129 (.A(b[18]), .ZN(n_1_930));
   INV_X1 i_1_1130 (.A(b[23]), .ZN(n_1_931));
   INV_X1 i_1_1131 (.A(b[25]), .ZN(n_1_932));
   INV_X1 i_1_1132 (.A(counter[0]), .ZN(n_1_933));
   INV_X1 i_1_1133 (.A(counter[1]), .ZN(n_1_934));
   INV_X1 i_1_1134 (.A(counter[2]), .ZN(n_1_935));
   INV_X1 i_1_1135 (.A(counter[3]), .ZN(n_1_936));
   INV_X1 i_1_1136 (.A(counter[4]), .ZN(n_1_937));
   AOI21_X1 i_1_1137 (.A(n_1_728), .B1(n_1_704), .B2(n_1_701), .ZN(n_1_938));
   CLKGATETST_X1 clk_gate_result_reg (.CK(clk), .E(n_266), .SE(1'b0), .GCK(n_0));
   DFF_X1 \result_reg[63]  (.D(n_131), .CK(n_0), .Q(result[63]), .QN());
   DFF_X1 \result_reg[62]  (.D(n_130), .CK(n_0), .Q(result[62]), .QN());
   DFF_X1 \result_reg[61]  (.D(n_129), .CK(n_0), .Q(result[61]), .QN());
   DFF_X1 \result_reg[60]  (.D(n_128), .CK(n_0), .Q(result[60]), .QN());
   DFF_X1 \result_reg[59]  (.D(n_127), .CK(n_0), .Q(result[59]), .QN());
   DFF_X1 \result_reg[58]  (.D(n_126), .CK(n_0), .Q(result[58]), .QN());
   DFF_X1 \result_reg[57]  (.D(n_125), .CK(n_0), .Q(result[57]), .QN());
   DFF_X1 \result_reg[56]  (.D(n_124), .CK(n_0), .Q(result[56]), .QN());
   DFF_X1 \result_reg[55]  (.D(n_123), .CK(n_0), .Q(result[55]), .QN());
   DFF_X1 \result_reg[54]  (.D(n_122), .CK(n_0), .Q(result[54]), .QN());
   DFF_X1 \result_reg[53]  (.D(n_121), .CK(n_0), .Q(result[53]), .QN());
   DFF_X1 \result_reg[52]  (.D(n_120), .CK(n_0), .Q(result[52]), .QN());
   DFF_X1 \result_reg[51]  (.D(n_119), .CK(n_0), .Q(result[51]), .QN());
   DFF_X1 \result_reg[50]  (.D(n_118), .CK(n_0), .Q(result[50]), .QN());
   DFF_X1 \result_reg[49]  (.D(n_117), .CK(n_0), .Q(result[49]), .QN());
   DFF_X1 \result_reg[48]  (.D(n_116), .CK(n_0), .Q(result[48]), .QN());
   DFF_X1 \result_reg[47]  (.D(n_115), .CK(n_0), .Q(result[47]), .QN());
   DFF_X1 \result_reg[46]  (.D(n_114), .CK(n_0), .Q(result[46]), .QN());
   DFF_X1 \result_reg[45]  (.D(n_113), .CK(n_0), .Q(result[45]), .QN());
   DFF_X1 \result_reg[44]  (.D(n_112), .CK(n_0), .Q(result[44]), .QN());
   DFF_X1 \result_reg[43]  (.D(n_111), .CK(n_0), .Q(result[43]), .QN());
   DFF_X1 \result_reg[42]  (.D(n_110), .CK(n_0), .Q(result[42]), .QN());
   DFF_X1 \result_reg[41]  (.D(n_109), .CK(n_0), .Q(result[41]), .QN());
   DFF_X1 \result_reg[40]  (.D(n_108), .CK(n_0), .Q(result[40]), .QN());
   DFF_X1 \result_reg[39]  (.D(n_107), .CK(n_0), .Q(result[39]), .QN());
   DFF_X1 \result_reg[38]  (.D(n_106), .CK(n_0), .Q(result[38]), .QN());
   DFF_X1 \result_reg[37]  (.D(n_105), .CK(n_0), .Q(result[37]), .QN());
   DFF_X1 \result_reg[36]  (.D(n_104), .CK(n_0), .Q(result[36]), .QN());
   DFF_X1 \result_reg[35]  (.D(n_103), .CK(n_0), .Q(result[35]), .QN());
   DFF_X1 \result_reg[34]  (.D(n_102), .CK(n_0), .Q(result[34]), .QN());
   DFF_X1 \result_reg[33]  (.D(n_101), .CK(n_0), .Q(result[33]), .QN());
   DFF_X1 \result_reg[32]  (.D(n_100), .CK(n_0), .Q(result[32]), .QN());
   DFF_X1 \result_reg[31]  (.D(n_99), .CK(n_0), .Q(result[31]), .QN());
   DFF_X1 \result_reg[30]  (.D(n_98), .CK(n_0), .Q(result[30]), .QN());
   DFF_X1 \result_reg[29]  (.D(n_97), .CK(n_0), .Q(result[29]), .QN());
   DFF_X1 \result_reg[28]  (.D(n_96), .CK(n_0), .Q(result[28]), .QN());
   DFF_X1 \result_reg[27]  (.D(n_95), .CK(n_0), .Q(result[27]), .QN());
   DFF_X1 \result_reg[26]  (.D(n_94), .CK(n_0), .Q(result[26]), .QN());
   DFF_X1 \result_reg[25]  (.D(n_93), .CK(n_0), .Q(result[25]), .QN());
   DFF_X1 \result_reg[24]  (.D(n_92), .CK(n_0), .Q(result[24]), .QN());
   DFF_X1 \result_reg[23]  (.D(n_91), .CK(n_0), .Q(result[23]), .QN());
   DFF_X1 \result_reg[22]  (.D(n_90), .CK(n_0), .Q(result[22]), .QN());
   DFF_X1 \result_reg[21]  (.D(n_89), .CK(n_0), .Q(result[21]), .QN());
   DFF_X1 \result_reg[20]  (.D(n_88), .CK(n_0), .Q(result[20]), .QN());
   DFF_X1 \result_reg[19]  (.D(n_87), .CK(n_0), .Q(result[19]), .QN());
   DFF_X1 \result_reg[18]  (.D(n_86), .CK(n_0), .Q(result[18]), .QN());
   DFF_X1 \result_reg[17]  (.D(n_85), .CK(n_0), .Q(result[17]), .QN());
   DFF_X1 \result_reg[16]  (.D(n_84), .CK(n_0), .Q(result[16]), .QN());
   DFF_X1 \result_reg[15]  (.D(n_83), .CK(n_0), .Q(result[15]), .QN());
   DFF_X1 \result_reg[14]  (.D(n_82), .CK(n_0), .Q(result[14]), .QN());
   DFF_X1 \result_reg[13]  (.D(n_81), .CK(n_0), .Q(result[13]), .QN());
   DFF_X1 \result_reg[12]  (.D(n_80), .CK(n_0), .Q(result[12]), .QN());
   DFF_X1 \result_reg[11]  (.D(n_79), .CK(n_0), .Q(result[11]), .QN());
   DFF_X1 \result_reg[10]  (.D(n_78), .CK(n_0), .Q(result[10]), .QN());
   DFF_X1 \result_reg[9]  (.D(n_77), .CK(n_0), .Q(result[9]), .QN());
   DFF_X1 \result_reg[8]  (.D(n_76), .CK(n_0), .Q(result[8]), .QN());
   DFF_X1 \result_reg[7]  (.D(n_75), .CK(n_0), .Q(result[7]), .QN());
   DFF_X1 \result_reg[6]  (.D(n_74), .CK(n_0), .Q(result[6]), .QN());
   DFF_X1 \result_reg[5]  (.D(n_73), .CK(n_0), .Q(result[5]), .QN());
   DFF_X1 \result_reg[4]  (.D(n_72), .CK(n_0), .Q(result[4]), .QN());
   DFF_X1 \result_reg[3]  (.D(n_71), .CK(n_0), .Q(result[3]), .QN());
   DFF_X1 \result_reg[2]  (.D(n_70), .CK(n_0), .Q(result[2]), .QN());
   DFF_X1 \result_reg[1]  (.D(n_69), .CK(n_0), .Q(result[1]), .QN());
   DFF_X1 \result_reg[0]  (.D(n_68), .CK(n_0), .Q(result[0]), .QN());
   CLKGATETST_X1 clk_gate_counter_reg (.CK(clk), .E(en), .SE(1'b0), .GCK(n_1));
   DFF_X1 \counter_reg[4]  (.D(n_136), .CK(n_1), .Q(counter[4]), .QN());
   DFF_X1 \counter_reg[3]  (.D(n_135), .CK(n_1), .Q(counter[3]), .QN());
   DFF_X1 \counter_reg[2]  (.D(n_134), .CK(n_1), .Q(counter[2]), .QN());
   DFF_X1 \counter_reg[1]  (.D(n_133), .CK(n_1), .Q(counter[1]), .QN());
   DFF_X1 \counter_reg[0]  (.D(n_132), .CK(n_1), .Q(counter[0]), .QN());
   DFF_X1 resetReg_reg (.D(n_269), .CK(clk), .Q(resetReg), .QN());
   MUX2_X1 resetReg_reg_enable_mux_0 (.A(resetReg), .B(n_67), .S(n_267), 
      .Z(n_269));
   CLKGATETST_X1 clk_gate_aux_reg (.CK(clk), .E(n_265), .SE(1'b0), .GCK(n_2));
   DFF_X1 \aux_reg[63]  (.D(n_200), .CK(n_2), .Q(aux[63]), .QN());
   DFF_X1 \aux_reg[62]  (.D(n_199), .CK(n_2), .Q(aux[62]), .QN());
   DFF_X1 \aux_reg[61]  (.D(n_198), .CK(n_2), .Q(aux[61]), .QN());
   DFF_X1 \aux_reg[60]  (.D(n_197), .CK(n_2), .Q(aux[60]), .QN());
   DFF_X1 \aux_reg[59]  (.D(n_196), .CK(n_2), .Q(aux[59]), .QN());
   DFF_X1 \aux_reg[58]  (.D(n_195), .CK(n_2), .Q(aux[58]), .QN());
   DFF_X1 \aux_reg[57]  (.D(n_194), .CK(n_2), .Q(aux[57]), .QN());
   DFF_X1 \aux_reg[56]  (.D(n_193), .CK(n_2), .Q(aux[56]), .QN());
   DFF_X1 \aux_reg[55]  (.D(n_192), .CK(n_2), .Q(aux[55]), .QN());
   DFF_X1 \aux_reg[54]  (.D(n_191), .CK(n_2), .Q(aux[54]), .QN());
   DFF_X1 \aux_reg[53]  (.D(n_190), .CK(n_2), .Q(aux[53]), .QN());
   DFF_X1 \aux_reg[52]  (.D(n_189), .CK(n_2), .Q(aux[52]), .QN());
   DFF_X1 \aux_reg[51]  (.D(n_188), .CK(n_2), .Q(aux[51]), .QN());
   DFF_X1 \aux_reg[50]  (.D(n_187), .CK(n_2), .Q(aux[50]), .QN());
   DFF_X1 \aux_reg[49]  (.D(n_186), .CK(n_2), .Q(aux[49]), .QN());
   DFF_X1 \aux_reg[48]  (.D(n_185), .CK(n_2), .Q(aux[48]), .QN());
   DFF_X1 \aux_reg[47]  (.D(n_184), .CK(n_2), .Q(aux[47]), .QN());
   DFF_X1 \aux_reg[46]  (.D(n_183), .CK(n_2), .Q(aux[46]), .QN());
   DFF_X1 \aux_reg[45]  (.D(n_182), .CK(n_2), .Q(aux[45]), .QN());
   DFF_X1 \aux_reg[44]  (.D(n_181), .CK(n_2), .Q(aux[44]), .QN());
   DFF_X1 \aux_reg[43]  (.D(n_180), .CK(n_2), .Q(aux[43]), .QN());
   DFF_X1 \aux_reg[42]  (.D(n_179), .CK(n_2), .Q(aux[42]), .QN());
   DFF_X1 \aux_reg[41]  (.D(n_178), .CK(n_2), .Q(aux[41]), .QN());
   DFF_X1 \aux_reg[40]  (.D(n_177), .CK(n_2), .Q(aux[40]), .QN());
   DFF_X1 \aux_reg[39]  (.D(n_176), .CK(n_2), .Q(aux[39]), .QN());
   DFF_X1 \aux_reg[38]  (.D(n_175), .CK(n_2), .Q(aux[38]), .QN());
   DFF_X1 \aux_reg[37]  (.D(n_174), .CK(n_2), .Q(aux[37]), .QN());
   DFF_X1 \aux_reg[36]  (.D(n_173), .CK(n_2), .Q(aux[36]), .QN());
   DFF_X1 \aux_reg[35]  (.D(n_172), .CK(n_2), .Q(aux[35]), .QN());
   DFF_X1 \aux_reg[34]  (.D(n_171), .CK(n_2), .Q(aux[34]), .QN());
   DFF_X1 \aux_reg[33]  (.D(n_170), .CK(n_2), .Q(aux[33]), .QN());
   DFF_X1 \aux_reg[32]  (.D(n_169), .CK(n_2), .Q(aux[32]), .QN());
   DFF_X1 \aux_reg[31]  (.D(n_168), .CK(n_2), .Q(aux[31]), .QN());
   DFF_X1 \aux_reg[30]  (.D(n_167), .CK(n_2), .Q(aux[30]), .QN());
   DFF_X1 \aux_reg[29]  (.D(n_166), .CK(n_2), .Q(aux[29]), .QN());
   DFF_X1 \aux_reg[28]  (.D(n_165), .CK(n_2), .Q(aux[28]), .QN());
   DFF_X1 \aux_reg[27]  (.D(n_164), .CK(n_2), .Q(aux[27]), .QN());
   DFF_X1 \aux_reg[26]  (.D(n_163), .CK(n_2), .Q(aux[26]), .QN());
   DFF_X1 \aux_reg[25]  (.D(n_162), .CK(n_2), .Q(aux[25]), .QN());
   DFF_X1 \aux_reg[24]  (.D(n_161), .CK(n_2), .Q(aux[24]), .QN());
   DFF_X1 \aux_reg[23]  (.D(n_160), .CK(n_2), .Q(aux[23]), .QN());
   DFF_X1 \aux_reg[22]  (.D(n_159), .CK(n_2), .Q(aux[22]), .QN());
   DFF_X1 \aux_reg[21]  (.D(n_158), .CK(n_2), .Q(aux[21]), .QN());
   DFF_X1 \aux_reg[20]  (.D(n_157), .CK(n_2), .Q(aux[20]), .QN());
   DFF_X1 \aux_reg[19]  (.D(n_156), .CK(n_2), .Q(aux[19]), .QN());
   DFF_X1 \aux_reg[18]  (.D(n_155), .CK(n_2), .Q(aux[18]), .QN());
   DFF_X1 \aux_reg[17]  (.D(n_154), .CK(n_2), .Q(aux[17]), .QN());
   DFF_X1 \aux_reg[16]  (.D(n_153), .CK(n_2), .Q(aux[16]), .QN());
   DFF_X1 \aux_reg[15]  (.D(n_152), .CK(n_2), .Q(aux[15]), .QN());
   DFF_X1 \aux_reg[14]  (.D(n_151), .CK(n_2), .Q(aux[14]), .QN());
   DFF_X1 \aux_reg[13]  (.D(n_150), .CK(n_2), .Q(aux[13]), .QN());
   DFF_X1 \aux_reg[12]  (.D(n_149), .CK(n_2), .Q(aux[12]), .QN());
   DFF_X1 \aux_reg[11]  (.D(n_148), .CK(n_2), .Q(aux[11]), .QN());
   DFF_X1 \aux_reg[10]  (.D(n_147), .CK(n_2), .Q(aux[10]), .QN());
   DFF_X1 \aux_reg[9]  (.D(n_146), .CK(n_2), .Q(aux[9]), .QN());
   DFF_X1 \aux_reg[8]  (.D(n_145), .CK(n_2), .Q(aux[8]), .QN());
   DFF_X1 \aux_reg[7]  (.D(n_144), .CK(n_2), .Q(aux[7]), .QN());
   DFF_X1 \aux_reg[6]  (.D(n_143), .CK(n_2), .Q(aux[6]), .QN());
   DFF_X1 \aux_reg[5]  (.D(n_142), .CK(n_2), .Q(aux[5]), .QN());
   DFF_X1 \aux_reg[4]  (.D(n_141), .CK(n_2), .Q(aux[4]), .QN());
   DFF_X1 \aux_reg[3]  (.D(n_140), .CK(n_2), .Q(aux[3]), .QN());
   DFF_X1 \aux_reg[2]  (.D(n_139), .CK(n_2), .Q(aux[2]), .QN());
   DFF_X1 \aux_reg[1]  (.D(n_138), .CK(n_2), .Q(aux[1]), .QN());
   DFF_X1 \aux_reg[0]  (.D(n_137), .CK(n_2), .Q(aux[0]), .QN());
endmodule

module registerNbits__0_90(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module integrationMult(inputA, inputB, clk, reset, en, result);
   input [31:0]inputA;
   input [31:0]inputB;
   input clk;
   input reset;
   input en;
   output [63:0]result;

   wire [31:0]A_reg;
   wire [31:0]B_reg;
   wire enableOutput;
   wire [31:0]outB_reg;
   wire [31:0]outA_reg;

   registerNbits__0_84 regA (.clk(clk), .reset(reset), .en(en), .inp(inputA), 
      .out(A_reg));
   registerNbits__0_87 regB (.clk(clk), .reset(reset), .en(en), .inp(inputB), 
      .out(B_reg));
   radix4Booth radix4BoothIns (.a(A_reg), .b(B_reg), .clk(clk), .reset(reset), 
      .en(en), .result({outA_reg[31], outA_reg[30], outA_reg[29], outA_reg[28], 
      outA_reg[27], outA_reg[26], outA_reg[25], outA_reg[24], outA_reg[23], 
      outA_reg[22], outA_reg[21], outA_reg[20], outA_reg[19], outA_reg[18], 
      outA_reg[17], outA_reg[16], outA_reg[15], outA_reg[14], outA_reg[13], 
      outA_reg[12], outA_reg[11], outA_reg[10], outA_reg[9], outA_reg[8], 
      outA_reg[7], outA_reg[6], outA_reg[5], outA_reg[4], outA_reg[3], 
      outA_reg[2], outA_reg[1], outA_reg[0], outB_reg[31], outB_reg[30], 
      outB_reg[29], outB_reg[28], outB_reg[27], outB_reg[26], outB_reg[25], 
      outB_reg[24], outB_reg[23], outB_reg[22], outB_reg[21], outB_reg[20], 
      outB_reg[19], outB_reg[18], outB_reg[17], outB_reg[16], outB_reg[15], 
      outB_reg[14], outB_reg[13], outB_reg[12], outB_reg[11], outB_reg[10], 
      outB_reg[9], outB_reg[8], outB_reg[7], outB_reg[6], outB_reg[5], 
      outB_reg[4], outB_reg[3], outB_reg[2], outB_reg[1], outB_reg[0]}), 
      .enableOutput(enableOutput));
   registerNbits__0_90 outB (.clk(clk), .reset(reset), .en(enableOutput), 
      .inp(outA_reg), .out({result[63], result[62], result[61], result[60], 
      result[59], result[58], result[57], result[56], result[55], result[54], 
      result[53], result[52], result[51], result[50], result[49], result[48], 
      result[47], result[46], result[45], result[44], result[43], result[42], 
      result[41], result[40], result[39], result[38], result[37], result[36], 
      result[35], result[34], result[33], result[32]}));
   registerNbits outA (.clk(clk), .reset(reset), .en(enableOutput), .inp(
      outB_reg), .out({result[31], result[30], result[29], result[28], 
      result[27], result[26], result[25], result[24], result[23], result[22], 
      result[21], result[20], result[19], result[18], result[17], result[16], 
      result[15], result[14], result[13], result[12], result[11], result[10], 
      result[9], result[8], result[7], result[6], result[5], result[4], 
      result[3], result[2], result[1], result[0]}));
endmodule
