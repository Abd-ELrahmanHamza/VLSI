
// 	Fri Dec 23 02:56:30 2022
//	vlsi
//	192.168.219.129

module registerNbits__parameterized0 (clk__CTS_1_PP_35, clk__CTS_1_PP_36, clk__CTS_1_PP_2, 
    clk__CTS_1_PP_3, clk__CTS_1_PP_41, clk, inp, out);

output [63:0] out;
output clk__CTS_1_PP_35;
output clk__CTS_1_PP_36;
input clk;
input [63:0] inp;
input clk__CTS_1_PP_2;
input clk__CTS_1_PP_3;
input clk__CTS_1_PP_41;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk__CTS_1_PP_3), .D (inp[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk__CTS_1_PP_3), .D (inp[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk__CTS_1_PP_3), .D (inp[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk__CTS_1_PP_3), .D (inp[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk__CTS_1_PP_3), .D (inp[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk__CTS_1_PP_3), .D (inp[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk__CTS_1_PP_3), .D (inp[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk__CTS_1_PP_3), .D (inp[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk__CTS_1_PP_3), .D (inp[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk__CTS_1_PP_3), .D (inp[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk__CTS_1_PP_3), .D (inp[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk__CTS_1_PP_3), .D (inp[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk__CTS_1_PP_3), .D (inp[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk__CTS_1_PP_3), .D (inp[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk__CTS_1_PP_3), .D (inp[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk__CTS_1_PP_3), .D (inp[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk__CTS_1_PP_3), .D (inp[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk__CTS_1_PP_36), .D (inp[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk__CTS_1_PP_36), .D (inp[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk__CTS_1_PP_36), .D (inp[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk__CTS_1_PP_36), .D (inp[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk__CTS_1_PP_36), .D (inp[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk__CTS_1_PP_36), .D (inp[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk__CTS_1_PP_36), .D (inp[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk__CTS_1_PP_36), .D (inp[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk__CTS_1_PP_36), .D (inp[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk__CTS_1_PP_36), .D (inp[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk__CTS_1_PP_36), .D (inp[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk__CTS_1_PP_36), .D (inp[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk__CTS_1_PP_36), .D (inp[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk__CTS_1_PP_36), .D (inp[30]));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk__CTS_1_PP_36), .D (inp[31]));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (clk__CTS_1_PP_3), .D (inp[32]));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (clk__CTS_1_PP_3), .D (inp[33]));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (clk__CTS_1_PP_36), .D (inp[34]));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (clk__CTS_1_PP_36), .D (inp[35]));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (clk__CTS_1_PP_36), .D (inp[36]));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (clk__CTS_1_PP_36), .D (inp[37]));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (clk__CTS_1_PP_36), .D (inp[38]));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (clk__CTS_1_PP_35), .D (inp[39]));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (clk__CTS_1_PP_35), .D (inp[40]));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (clk__CTS_1_PP_35), .D (inp[41]));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (clk__CTS_1_PP_35), .D (inp[42]));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (clk__CTS_1_PP_35), .D (inp[43]));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (clk__CTS_1_PP_35), .D (inp[44]));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (clk__CTS_1_PP_35), .D (inp[45]));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (clk__CTS_1_PP_35), .D (inp[46]));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (clk__CTS_1_PP_35), .D (inp[47]));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (clk__CTS_1_PP_35), .D (inp[48]));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (clk__CTS_1_PP_2), .D (inp[49]));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (clk__CTS_1_PP_2), .D (inp[50]));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (clk__CTS_1_PP_2), .D (inp[51]));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (clk__CTS_1_PP_2), .D (inp[52]));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (clk__CTS_1_PP_2), .D (inp[53]));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (clk__CTS_1_PP_2), .D (inp[54]));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (clk__CTS_1_PP_2), .D (inp[55]));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (clk__CTS_1_PP_2), .D (inp[56]));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (clk__CTS_1_PP_2), .D (inp[57]));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (clk__CTS_1_PP_3), .D (inp[58]));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (clk__CTS_1_PP_3), .D (inp[59]));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (clk__CTS_1_PP_3), .D (inp[60]));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (clk__CTS_1_PP_2), .D (inp[61]));
DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (clk__CTS_1_PP_2), .D (inp[63]));
INV_X4 CTS_L9_c_tid1_9 (.ZN (clk__CTS_1_PP_35), .A (clk__CTS_1_PP_41));
INV_X4 CTS_L9_c_tid1_10 (.ZN (clk__CTS_1_PP_36), .A (clk__CTS_1_PP_41));

endmodule //registerNbits__parameterized0

module datapath__0_31 (a, p_0, m);

output [31:0] p_0;
input [31:0] a;
input [31:0] m;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;


XNOR2_X1 i_126 (.ZN (p_0[31]), .A (n_94), .B (m[31]));
OAI33_X1 i_125 (.ZN (n_94), .A1 (n_93), .A2 (a[31]), .A3 (m[30]), .B1 (n_89), .B2 (n_90), .B3 (n_91));
INV_X1 i_124 (.ZN (n_93), .A (n_89));
XNOR2_X1 i_123 (.ZN (p_0[30]), .A (n_89), .B (n_92));
AOI22_X1 i_122 (.ZN (n_92), .A1 (n_90), .A2 (n_91), .B1 (a[31]), .B2 (m[30]));
INV_X1 i_121 (.ZN (n_91), .A (m[30]));
INV_X1 i_120 (.ZN (n_90), .A (a[31]));
AOI22_X1 i_119 (.ZN (n_89), .A1 (n_86), .A2 (n_87), .B1 (n_88), .B2 (m[29]));
INV_X1 i_118 (.ZN (n_88), .A (a[29]));
XNOR2_X1 i_117 (.ZN (p_0[29]), .A (n_86), .B (n_87));
XNOR2_X1 i_116 (.ZN (n_87), .A (a[29]), .B (m[29]));
OAI22_X1 i_115 (.ZN (n_86), .A1 (n_83), .A2 (n_84), .B1 (n_85), .B2 (a[28]));
INV_X1 i_114 (.ZN (n_85), .A (m[28]));
XNOR2_X1 i_113 (.ZN (p_0[28]), .A (n_83), .B (n_84));
XOR2_X1 i_112 (.Z (n_84), .A (a[28]), .B (m[28]));
AOI22_X1 i_111 (.ZN (n_83), .A1 (n_80), .A2 (n_81), .B1 (n_82), .B2 (m[27]));
INV_X1 i_110 (.ZN (n_82), .A (a[27]));
XNOR2_X1 i_109 (.ZN (p_0[27]), .A (n_80), .B (n_81));
XNOR2_X1 i_108 (.ZN (n_81), .A (a[27]), .B (m[27]));
OAI22_X1 i_107 (.ZN (n_80), .A1 (n_77), .A2 (n_78), .B1 (n_79), .B2 (a[26]));
INV_X1 i_106 (.ZN (n_79), .A (m[26]));
XNOR2_X1 i_105 (.ZN (p_0[26]), .A (n_77), .B (n_78));
XOR2_X1 i_104 (.Z (n_78), .A (a[26]), .B (m[26]));
AOI22_X1 i_103 (.ZN (n_77), .A1 (n_74), .A2 (n_75), .B1 (n_76), .B2 (m[25]));
INV_X1 i_102 (.ZN (n_76), .A (a[25]));
XNOR2_X1 i_101 (.ZN (p_0[25]), .A (n_74), .B (n_75));
XNOR2_X1 i_100 (.ZN (n_75), .A (a[25]), .B (m[25]));
OAI22_X1 i_99 (.ZN (n_74), .A1 (n_71), .A2 (n_72), .B1 (n_73), .B2 (a[24]));
INV_X1 i_98 (.ZN (n_73), .A (m[24]));
XNOR2_X1 i_97 (.ZN (p_0[24]), .A (n_71), .B (n_72));
XOR2_X1 i_96 (.Z (n_72), .A (a[24]), .B (m[24]));
AOI22_X1 i_95 (.ZN (n_71), .A1 (n_68), .A2 (n_69), .B1 (n_70), .B2 (m[23]));
INV_X1 i_94 (.ZN (n_70), .A (a[23]));
XNOR2_X1 i_93 (.ZN (p_0[23]), .A (n_68), .B (n_69));
XNOR2_X1 i_92 (.ZN (n_69), .A (a[23]), .B (m[23]));
OAI22_X1 i_91 (.ZN (n_68), .A1 (n_65), .A2 (n_66), .B1 (n_67), .B2 (a[22]));
INV_X1 i_90 (.ZN (n_67), .A (m[22]));
XNOR2_X1 i_89 (.ZN (p_0[22]), .A (n_65), .B (n_66));
XOR2_X1 i_88 (.Z (n_66), .A (a[22]), .B (m[22]));
AOI22_X1 i_87 (.ZN (n_65), .A1 (n_62), .A2 (n_63), .B1 (n_64), .B2 (m[21]));
INV_X1 i_86 (.ZN (n_64), .A (a[21]));
XNOR2_X1 i_85 (.ZN (p_0[21]), .A (n_62), .B (n_63));
XNOR2_X1 i_84 (.ZN (n_63), .A (a[21]), .B (m[21]));
OAI22_X1 i_83 (.ZN (n_62), .A1 (n_59), .A2 (n_60), .B1 (n_61), .B2 (a[20]));
INV_X1 i_82 (.ZN (n_61), .A (m[20]));
XNOR2_X1 i_81 (.ZN (p_0[20]), .A (n_59), .B (n_60));
XOR2_X1 i_80 (.Z (n_60), .A (a[20]), .B (m[20]));
AOI22_X1 i_79 (.ZN (n_59), .A1 (n_56), .A2 (n_57), .B1 (n_58), .B2 (m[19]));
INV_X1 i_78 (.ZN (n_58), .A (a[19]));
XNOR2_X1 i_77 (.ZN (p_0[19]), .A (n_56), .B (n_57));
XNOR2_X1 i_76 (.ZN (n_57), .A (a[19]), .B (m[19]));
OAI22_X1 i_75 (.ZN (n_56), .A1 (n_53), .A2 (n_54), .B1 (n_55), .B2 (a[18]));
INV_X1 i_74 (.ZN (n_55), .A (m[18]));
XNOR2_X1 i_73 (.ZN (p_0[18]), .A (n_53), .B (n_54));
XOR2_X1 i_72 (.Z (n_54), .A (a[18]), .B (m[18]));
AOI22_X1 i_71 (.ZN (n_53), .A1 (n_50), .A2 (n_51), .B1 (n_52), .B2 (m[17]));
INV_X1 i_70 (.ZN (n_52), .A (a[17]));
XNOR2_X1 i_69 (.ZN (p_0[17]), .A (n_50), .B (n_51));
XNOR2_X1 i_68 (.ZN (n_51), .A (a[17]), .B (m[17]));
OAI22_X1 i_67 (.ZN (n_50), .A1 (n_47), .A2 (n_48), .B1 (n_49), .B2 (a[16]));
INV_X1 i_66 (.ZN (n_49), .A (m[16]));
XNOR2_X1 i_65 (.ZN (p_0[16]), .A (n_47), .B (n_48));
XOR2_X1 i_64 (.Z (n_48), .A (a[16]), .B (m[16]));
AOI22_X1 i_63 (.ZN (n_47), .A1 (n_44), .A2 (n_45), .B1 (n_46), .B2 (m[15]));
INV_X1 i_62 (.ZN (n_46), .A (a[15]));
XNOR2_X1 i_61 (.ZN (p_0[15]), .A (n_44), .B (n_45));
XNOR2_X1 i_60 (.ZN (n_45), .A (a[15]), .B (m[15]));
OAI22_X1 i_59 (.ZN (n_44), .A1 (n_41), .A2 (n_42), .B1 (n_43), .B2 (a[14]));
INV_X1 i_58 (.ZN (n_43), .A (m[14]));
XNOR2_X1 i_57 (.ZN (p_0[14]), .A (n_41), .B (n_42));
XOR2_X1 i_56 (.Z (n_42), .A (a[14]), .B (m[14]));
AOI22_X1 i_55 (.ZN (n_41), .A1 (n_38), .A2 (n_39), .B1 (n_40), .B2 (m[13]));
INV_X1 i_54 (.ZN (n_40), .A (a[13]));
XNOR2_X1 i_53 (.ZN (p_0[13]), .A (n_38), .B (n_39));
XNOR2_X1 i_52 (.ZN (n_39), .A (a[13]), .B (m[13]));
OAI22_X1 i_51 (.ZN (n_38), .A1 (n_35), .A2 (n_36), .B1 (n_37), .B2 (a[12]));
INV_X1 i_50 (.ZN (n_37), .A (m[12]));
XNOR2_X1 i_49 (.ZN (p_0[12]), .A (n_35), .B (n_36));
XOR2_X1 i_48 (.Z (n_36), .A (a[12]), .B (m[12]));
AOI22_X1 i_47 (.ZN (n_35), .A1 (n_32), .A2 (n_33), .B1 (n_34), .B2 (m[11]));
INV_X1 i_46 (.ZN (n_34), .A (a[11]));
XNOR2_X1 i_45 (.ZN (p_0[11]), .A (n_32), .B (n_33));
XNOR2_X1 i_44 (.ZN (n_33), .A (a[11]), .B (m[11]));
OAI22_X1 i_43 (.ZN (n_32), .A1 (n_29), .A2 (n_30), .B1 (n_31), .B2 (a[10]));
INV_X1 i_42 (.ZN (n_31), .A (m[10]));
XNOR2_X1 i_41 (.ZN (p_0[10]), .A (n_29), .B (n_30));
XOR2_X1 i_40 (.Z (n_30), .A (a[10]), .B (m[10]));
AOI22_X1 i_39 (.ZN (n_29), .A1 (n_26), .A2 (n_27), .B1 (n_28), .B2 (m[9]));
INV_X1 i_38 (.ZN (n_28), .A (a[9]));
XNOR2_X1 i_37 (.ZN (p_0[9]), .A (n_26), .B (n_27));
XNOR2_X1 i_36 (.ZN (n_27), .A (a[9]), .B (m[9]));
OAI22_X1 i_35 (.ZN (n_26), .A1 (n_23), .A2 (n_24), .B1 (n_25), .B2 (a[8]));
INV_X1 i_34 (.ZN (n_25), .A (m[8]));
XNOR2_X1 i_33 (.ZN (p_0[8]), .A (n_23), .B (n_24));
XOR2_X1 i_32 (.Z (n_24), .A (a[8]), .B (m[8]));
AOI22_X1 i_31 (.ZN (n_23), .A1 (n_20), .A2 (n_21), .B1 (n_22), .B2 (m[7]));
INV_X1 i_30 (.ZN (n_22), .A (a[7]));
XNOR2_X1 i_29 (.ZN (p_0[7]), .A (n_20), .B (n_21));
XNOR2_X1 i_28 (.ZN (n_21), .A (a[7]), .B (m[7]));
OAI22_X1 i_27 (.ZN (n_20), .A1 (n_17), .A2 (n_18), .B1 (n_19), .B2 (a[6]));
INV_X1 i_26 (.ZN (n_19), .A (m[6]));
XNOR2_X1 i_25 (.ZN (p_0[6]), .A (n_17), .B (n_18));
XOR2_X1 i_24 (.Z (n_18), .A (a[6]), .B (m[6]));
AOI22_X1 i_23 (.ZN (n_17), .A1 (n_14), .A2 (n_15), .B1 (n_16), .B2 (m[5]));
INV_X1 i_22 (.ZN (n_16), .A (a[5]));
XNOR2_X1 i_21 (.ZN (p_0[5]), .A (n_14), .B (n_15));
XNOR2_X1 i_20 (.ZN (n_15), .A (a[5]), .B (m[5]));
OAI22_X1 i_19 (.ZN (n_14), .A1 (n_11), .A2 (n_12), .B1 (n_13), .B2 (a[4]));
INV_X1 i_18 (.ZN (n_13), .A (m[4]));
XNOR2_X1 i_17 (.ZN (p_0[4]), .A (n_11), .B (n_12));
XOR2_X1 i_16 (.Z (n_12), .A (a[4]), .B (m[4]));
AOI22_X1 i_15 (.ZN (n_11), .A1 (n_8), .A2 (n_9), .B1 (n_10), .B2 (m[3]));
INV_X1 i_14 (.ZN (n_10), .A (a[3]));
XNOR2_X1 i_13 (.ZN (p_0[3]), .A (n_8), .B (n_9));
XNOR2_X1 i_12 (.ZN (n_9), .A (a[3]), .B (m[3]));
OAI22_X1 i_11 (.ZN (n_8), .A1 (n_5), .A2 (n_6), .B1 (n_7), .B2 (a[2]));
INV_X1 i_10 (.ZN (n_7), .A (m[2]));
XNOR2_X1 i_9 (.ZN (p_0[2]), .A (n_5), .B (n_6));
XOR2_X1 i_8 (.Z (n_6), .A (m[2]), .B (a[2]));
AOI22_X1 i_7 (.ZN (n_5), .A1 (n_2), .A2 (n_3), .B1 (n_4), .B2 (m[1]));
INV_X1 i_6 (.ZN (n_4), .A (a[1]));
INV_X1 i_5 (.ZN (n_3), .A (n_1));
XOR2_X1 i_4 (.Z (p_0[1]), .A (n_2), .B (n_1));
XNOR2_X1 i_3 (.ZN (n_2), .A (a[1]), .B (m[1]));
OAI21_X1 i_2 (.ZN (p_0[0]), .A (n_1), .B1 (m[0]), .B2 (n_0));
NAND2_X1 i_1 (.ZN (n_1), .A1 (n_0), .A2 (m[0]));
INV_X1 i_0 (.ZN (n_0), .A (a[0]));

endmodule //datapath__0_31

module datapath (m, a, p_0);

output [31:0] p_0;
input [31:0] a;
input [31:0] m;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;


XNOR2_X1 i_32 (.ZN (p_0[31]), .A (n_31), .B (n_30));
XNOR2_X1 i_31 (.ZN (n_31), .A (m[31]), .B (a[31]));
FA_X1 i_30 (.CO (n_30), .S (p_0[30]), .A (m[30]), .B (a[31]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_0[29]), .A (m[29]), .B (a[29]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_0[28]), .A (m[28]), .B (a[28]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_0[27]), .A (m[27]), .B (a[27]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_0[26]), .A (m[26]), .B (a[26]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_0[25]), .A (m[25]), .B (a[25]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_0[24]), .A (m[24]), .B (a[24]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_0[23]), .A (m[23]), .B (a[23]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_0[22]), .A (m[22]), .B (a[22]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_0[21]), .A (m[21]), .B (a[21]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_0[20]), .A (m[20]), .B (a[20]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_0[19]), .A (m[19]), .B (a[19]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_0[18]), .A (m[18]), .B (a[18]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_0[17]), .A (m[17]), .B (a[17]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_0[16]), .A (m[16]), .B (a[16]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_0[15]), .A (m[15]), .B (a[15]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_0[14]), .A (m[14]), .B (a[14]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_0[13]), .A (m[13]), .B (a[13]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_0[12]), .A (m[12]), .B (a[12]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_0[11]), .A (m[11]), .B (a[11]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_0[10]), .A (m[10]), .B (a[10]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_0[9]), .A (m[9]), .B (a[9]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_0[8]), .A (m[8]), .B (a[8]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_0[7]), .A (m[7]), .B (a[7]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_0[6]), .A (m[6]), .B (a[6]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_0[5]), .A (m[5]), .B (a[5]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_0[4]), .A (m[4]), .B (a[4]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_0[3]), .A (m[3]), .B (a[3]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_0[2]), .A (m[2]), .B (a[2]), .CI (n_1));
FA_X1 i_1 (.CO (n_1), .S (p_0[1]), .A (m[1]), .B (a[1]), .CI (n_0));
HA_X1 i_0 (.CO (n_0), .S (p_0[0]), .A (m[0]), .B (a[0]));

endmodule //datapath

module booth_multiplier (clk__CTS_1_PP_0, clk__CTS_1_PP_1, in1, in2, clk, rst, out);

output [63:0] out;
output clk__CTS_1_PP_0;
input clk;
input [31:0] in1;
input [31:0] in2;
input rst;
input clk__CTS_1_PP_1;
wire CTS_n_tid1_14;
wire CLOCK_slh_n74;
wire n_2_0;
wire n_2_1;
wire n_2_2;
wire n_2_3;
wire n_2_4;
wire n_2_5;
wire n_2_6;
wire n_2_7;
wire n_2_8;
wire n_2_9;
wire n_2_10;
wire n_2_11;
wire n_2_12;
wire n_2_13;
wire n_2_14;
wire n_2_15;
wire n_2_16;
wire n_2_17;
wire n_2_18;
wire n_2_19;
wire n_2_20;
wire n_2_21;
wire n_2_22;
wire n_2_23;
wire n_2_24;
wire n_2_25;
wire n_2_26;
wire n_2_27;
wire n_2_28;
wire n_2_29;
wire n_2_30;
wire n_2_31;
wire n_2_32;
wire n_2_33;
wire n_2_34;
wire n_2_35;
wire n_2_36;
wire n_2_37;
wire n_2_38;
wire n_2_39;
wire \m[31] ;
wire \m[30] ;
wire \m[29] ;
wire \m[28] ;
wire \m[27] ;
wire \m[26] ;
wire \m[25] ;
wire \m[24] ;
wire \m[23] ;
wire \m[22] ;
wire \m[21] ;
wire \m[20] ;
wire \m[19] ;
wire \m[18] ;
wire \m[17] ;
wire \m[16] ;
wire \m[15] ;
wire \m[14] ;
wire \m[13] ;
wire \m[12] ;
wire \m[11] ;
wire \m[10] ;
wire \m[9] ;
wire \m[8] ;
wire \m[7] ;
wire \m[6] ;
wire \m[5] ;
wire \m[4] ;
wire \m[3] ;
wire \m[2] ;
wire \m[1] ;
wire \m[0] ;
wire q0;
wire uc_0;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire n_0;
wire uc_1;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_98;
wire drc_ipo_n6;
wire drc_ipo_n5;
wire CTS_n_tid1_29;
wire CTS_n_tid1_26;
wire CTS_n_tid1_30;


DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (CTS_n_tid1_14), .D (n_127));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_14), .D (n_64));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (CTS_n_tid1_14), .D (n_126));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (CTS_n_tid1_14), .D (n_125));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (CTS_n_tid1_14), .D (n_124));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (CTS_n_tid1_14), .D (n_123));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (CTS_n_tid1_14), .D (n_122));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (CTS_n_tid1_14), .D (n_121));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (CTS_n_tid1_14), .D (n_120));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (CTS_n_tid1_14), .D (n_119));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (CTS_n_tid1_14), .D (n_118));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (CTS_n_tid1_14), .D (n_117));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (CTS_n_tid1_14), .D (n_116));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (CTS_n_tid1_14), .D (n_115));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (CTS_n_tid1_14), .D (n_114));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (CTS_n_tid1_14), .D (n_113));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (CTS_n_tid1_14), .D (n_112));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (CTS_n_tid1_14), .D (n_111));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (CTS_n_tid1_14), .D (n_110));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (CTS_n_tid1_14), .D (n_109));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (CTS_n_tid1_14), .D (n_108));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (CTS_n_tid1_14), .D (n_107));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (CTS_n_tid1_14), .D (n_106));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (CTS_n_tid1_14), .D (n_105));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (CTS_n_tid1_14), .D (n_104));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (CTS_n_tid1_14), .D (n_103));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (CTS_n_tid1_14), .D (n_102));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (CTS_n_tid1_14), .D (n_101));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (CTS_n_tid1_14), .D (n_100));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (CTS_n_tid1_14), .D (n_99));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (CTS_n_tid1_14), .D (n_97));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (CTS_n_tid1_14), .D (n_96));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid1_14), .D (n_95));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_14), .D (n_94));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_14), .D (n_93));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_14), .D (n_92));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_14), .D (n_91));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_14), .D (n_90));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_14), .D (n_89));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_14), .D (n_88));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_14), .D (n_87));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_14), .D (n_86));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_14), .D (n_85));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_14), .D (n_84));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_14), .D (n_83));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_14), .D (n_82));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_14), .D (n_81));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_14), .D (n_80));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_14), .D (n_79));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_14), .D (n_78));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_14), .D (n_77));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_14), .D (n_76));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_14), .D (n_75));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_14), .D (n_74));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_14), .D (n_73));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_14), .D (n_72));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_14), .D (n_71));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_14), .D (n_70));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_14), .D (n_69));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_14), .D (n_68));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_14), .D (n_67));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_14), .D (n_66));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_14), .D (n_65));
DFF_X1 q0_reg (.Q (q0), .CK (CTS_n_tid1_14), .D (n_128));
DFF_X1 \m_reg[0]  (.Q (\m[0] ), .CK (n_98), .D (in1[0]));
DFF_X1 \m_reg[1]  (.Q (\m[1] ), .CK (n_98), .D (in1[1]));
DFF_X1 \m_reg[2]  (.Q (\m[2] ), .CK (n_98), .D (in1[2]));
DFF_X1 \m_reg[3]  (.Q (\m[3] ), .CK (n_98), .D (in1[3]));
DFF_X1 \m_reg[4]  (.Q (\m[4] ), .CK (n_98), .D (in1[4]));
DFF_X1 \m_reg[5]  (.Q (\m[5] ), .CK (n_98), .D (in1[5]));
DFF_X1 \m_reg[6]  (.Q (\m[6] ), .CK (n_98), .D (in1[6]));
DFF_X1 \m_reg[7]  (.Q (\m[7] ), .CK (n_98), .D (in1[7]));
DFF_X1 \m_reg[8]  (.Q (\m[8] ), .CK (n_98), .D (in1[8]));
DFF_X1 \m_reg[9]  (.Q (\m[9] ), .CK (n_98), .D (in1[9]));
DFF_X1 \m_reg[10]  (.Q (\m[10] ), .CK (n_98), .D (in1[10]));
DFF_X1 \m_reg[11]  (.Q (\m[11] ), .CK (n_98), .D (in1[11]));
DFF_X1 \m_reg[12]  (.Q (\m[12] ), .CK (n_98), .D (in1[12]));
DFF_X1 \m_reg[13]  (.Q (\m[13] ), .CK (n_98), .D (in1[13]));
DFF_X1 \m_reg[14]  (.Q (\m[14] ), .CK (n_98), .D (in1[14]));
DFF_X1 \m_reg[15]  (.Q (\m[15] ), .CK (n_98), .D (in1[15]));
DFF_X1 \m_reg[16]  (.Q (\m[16] ), .CK (n_98), .D (in1[16]));
DFF_X1 \m_reg[17]  (.Q (\m[17] ), .CK (n_98), .D (in1[17]));
DFF_X1 \m_reg[18]  (.Q (\m[18] ), .CK (n_98), .D (in1[18]));
DFF_X1 \m_reg[19]  (.Q (\m[19] ), .CK (n_98), .D (in1[19]));
DFF_X1 \m_reg[20]  (.Q (\m[20] ), .CK (n_98), .D (in1[20]));
DFF_X1 \m_reg[21]  (.Q (\m[21] ), .CK (n_98), .D (in1[21]));
DFF_X1 \m_reg[22]  (.Q (\m[22] ), .CK (n_98), .D (in1[22]));
DFF_X1 \m_reg[23]  (.Q (\m[23] ), .CK (n_98), .D (in1[23]));
DFF_X1 \m_reg[24]  (.Q (\m[24] ), .CK (n_98), .D (in1[24]));
DFF_X1 \m_reg[25]  (.Q (\m[25] ), .CK (n_98), .D (in1[25]));
DFF_X1 \m_reg[26]  (.Q (\m[26] ), .CK (n_98), .D (in1[26]));
DFF_X1 \m_reg[27]  (.Q (\m[27] ), .CK (n_98), .D (in1[27]));
DFF_X1 \m_reg[28]  (.Q (\m[28] ), .CK (n_98), .D (in1[28]));
DFF_X1 \m_reg[29]  (.Q (\m[29] ), .CK (n_98), .D (in1[29]));
DFF_X1 \m_reg[30]  (.Q (\m[30] ), .CK (n_98), .D (in1[30]));
DFF_X1 \m_reg[31]  (.Q (\m[31] ), .CK (n_98), .D (in1[31]));
CLKGATETST_X1 clk_gate_m_reg (.GCK (n_98), .CK (CTS_n_tid1_29), .E (rst), .SE (1'b0 ));
INV_X1 i_2_103 (.ZN (n_2_39), .A (out[0]));
INV_X1 i_2_102 (.ZN (n_2_38), .A (q0));
XNOR2_X1 i_2_101 (.ZN (n_2_37), .A (n_2_39), .B (q0));
NOR2_X4 i_2_100 (.ZN (n_2_36), .A1 (n_2_37), .A2 (CLOCK_slh_n74));
NAND2_X1 i_2_99 (.ZN (n_2_35), .A1 (out[63]), .A2 (n_2_36));
NOR2_X1 i_2_98 (.ZN (n_128), .A1 (n_2_39), .A2 (CLOCK_slh_n74));
NOR3_X1 i_2_97 (.ZN (n_2_34), .A1 (n_2_39), .A2 (q0), .A3 (rst));
NOR3_X1 i_2_96 (.ZN (n_2_33), .A1 (n_2_38), .A2 (rst), .A3 (out[0]));
AOI22_X1 i_2_95 (.ZN (n_2_32), .A1 (n_63), .A2 (drc_ipo_n5), .B1 (drc_ipo_n6), .B2 (n_31));
NAND2_X1 i_2_94 (.ZN (n_127), .A1 (n_2_35), .A2 (n_2_32));
AOI22_X1 i_2_93 (.ZN (n_2_31), .A1 (n_62), .A2 (drc_ipo_n5), .B1 (drc_ipo_n6), .B2 (n_30));
NAND2_X1 i_2_92 (.ZN (n_126), .A1 (n_2_35), .A2 (n_2_31));
AOI222_X1 i_2_91 (.ZN (n_2_30), .A1 (out[61]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_61)
    , .C1 (drc_ipo_n6), .C2 (n_29));
INV_X1 i_2_90 (.ZN (n_125), .A (n_2_30));
AOI222_X1 i_2_89 (.ZN (n_2_29), .A1 (out[60]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_60)
    , .C1 (drc_ipo_n6), .C2 (n_28));
INV_X1 i_2_88 (.ZN (n_124), .A (n_2_29));
AOI222_X1 i_2_87 (.ZN (n_2_28), .A1 (out[59]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_59)
    , .C1 (drc_ipo_n6), .C2 (n_27));
INV_X1 i_2_86 (.ZN (n_123), .A (n_2_28));
AOI222_X1 i_2_85 (.ZN (n_2_27), .A1 (out[58]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_58)
    , .C1 (drc_ipo_n6), .C2 (n_26));
INV_X1 i_2_84 (.ZN (n_122), .A (n_2_27));
AOI222_X1 i_2_83 (.ZN (n_2_26), .A1 (out[57]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_57)
    , .C1 (drc_ipo_n6), .C2 (n_25));
INV_X1 i_2_82 (.ZN (n_121), .A (n_2_26));
AOI222_X1 i_2_81 (.ZN (n_2_25), .A1 (out[56]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_56)
    , .C1 (drc_ipo_n6), .C2 (n_24));
INV_X1 i_2_80 (.ZN (n_120), .A (n_2_25));
AOI222_X1 i_2_79 (.ZN (n_2_24), .A1 (out[55]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_55)
    , .C1 (drc_ipo_n6), .C2 (n_23));
INV_X1 i_2_78 (.ZN (n_119), .A (n_2_24));
AOI222_X1 i_2_77 (.ZN (n_2_23), .A1 (out[54]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_54)
    , .C1 (drc_ipo_n6), .C2 (n_22));
INV_X1 i_2_76 (.ZN (n_118), .A (n_2_23));
AOI222_X1 i_2_75 (.ZN (n_2_22), .A1 (out[53]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_53)
    , .C1 (drc_ipo_n6), .C2 (n_21));
INV_X1 i_2_74 (.ZN (n_117), .A (n_2_22));
AOI222_X1 i_2_73 (.ZN (n_2_21), .A1 (out[52]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_52)
    , .C1 (drc_ipo_n6), .C2 (n_20));
INV_X1 i_2_72 (.ZN (n_116), .A (n_2_21));
AOI222_X1 i_2_71 (.ZN (n_2_20), .A1 (out[51]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_51)
    , .C1 (drc_ipo_n6), .C2 (n_19));
INV_X1 i_2_70 (.ZN (n_115), .A (n_2_20));
AOI222_X1 i_2_69 (.ZN (n_2_19), .A1 (out[50]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_50)
    , .C1 (drc_ipo_n6), .C2 (n_18));
INV_X1 i_2_68 (.ZN (n_114), .A (n_2_19));
AOI222_X1 i_2_67 (.ZN (n_2_18), .A1 (out[49]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_49)
    , .C1 (drc_ipo_n6), .C2 (n_17));
INV_X1 i_2_66 (.ZN (n_113), .A (n_2_18));
AOI222_X1 i_2_65 (.ZN (n_2_17), .A1 (out[48]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_48)
    , .C1 (drc_ipo_n6), .C2 (n_16));
INV_X1 i_2_64 (.ZN (n_112), .A (n_2_17));
AOI222_X1 i_2_63 (.ZN (n_2_16), .A1 (out[47]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_47)
    , .C1 (drc_ipo_n6), .C2 (n_15));
INV_X1 i_2_62 (.ZN (n_111), .A (n_2_16));
AOI222_X1 i_2_61 (.ZN (n_2_15), .A1 (out[46]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_46)
    , .C1 (drc_ipo_n6), .C2 (n_14));
INV_X1 i_2_60 (.ZN (n_110), .A (n_2_15));
AOI222_X1 i_2_59 (.ZN (n_2_14), .A1 (out[45]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_45)
    , .C1 (drc_ipo_n6), .C2 (n_13));
INV_X1 i_2_58 (.ZN (n_109), .A (n_2_14));
AOI222_X1 i_2_57 (.ZN (n_2_13), .A1 (out[44]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_44)
    , .C1 (drc_ipo_n6), .C2 (n_12));
INV_X1 i_2_56 (.ZN (n_108), .A (n_2_13));
AOI222_X1 i_2_55 (.ZN (n_2_12), .A1 (out[43]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_43)
    , .C1 (drc_ipo_n6), .C2 (n_11));
INV_X1 i_2_54 (.ZN (n_107), .A (n_2_12));
AOI222_X1 i_2_53 (.ZN (n_2_11), .A1 (out[42]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_42)
    , .C1 (drc_ipo_n6), .C2 (n_10));
INV_X1 i_2_52 (.ZN (n_106), .A (n_2_11));
AOI222_X1 i_2_51 (.ZN (n_2_10), .A1 (out[41]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_41)
    , .C1 (drc_ipo_n6), .C2 (n_9));
INV_X1 i_2_50 (.ZN (n_105), .A (n_2_10));
AOI222_X1 i_2_49 (.ZN (n_2_9), .A1 (out[40]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_40)
    , .C1 (drc_ipo_n6), .C2 (n_8));
INV_X1 i_2_48 (.ZN (n_104), .A (n_2_9));
AOI222_X1 i_2_47 (.ZN (n_2_8), .A1 (out[39]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_39)
    , .C1 (drc_ipo_n6), .C2 (n_7));
INV_X1 i_2_46 (.ZN (n_103), .A (n_2_8));
AOI222_X1 i_2_45 (.ZN (n_2_7), .A1 (out[38]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_38)
    , .C1 (drc_ipo_n6), .C2 (n_6));
INV_X1 i_2_44 (.ZN (n_102), .A (n_2_7));
AOI222_X1 i_2_43 (.ZN (n_2_6), .A1 (out[37]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_37)
    , .C1 (drc_ipo_n6), .C2 (n_5));
INV_X1 i_2_42 (.ZN (n_101), .A (n_2_6));
AOI222_X1 i_2_41 (.ZN (n_2_5), .A1 (out[36]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_36)
    , .C1 (drc_ipo_n6), .C2 (n_4));
INV_X1 i_2_40 (.ZN (n_100), .A (n_2_5));
AOI222_X1 i_2_39 (.ZN (n_2_4), .A1 (out[35]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_35)
    , .C1 (drc_ipo_n6), .C2 (n_3));
INV_X1 i_2_38 (.ZN (n_99), .A (n_2_4));
AOI222_X1 i_2_37 (.ZN (n_2_3), .A1 (out[34]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_34)
    , .C1 (drc_ipo_n6), .C2 (n_2));
INV_X1 i_2_36 (.ZN (n_97), .A (n_2_3));
AOI222_X1 i_2_35 (.ZN (n_2_2), .A1 (out[33]), .A2 (n_2_36), .B1 (drc_ipo_n5), .B2 (n_33)
    , .C1 (drc_ipo_n6), .C2 (n_1));
INV_X1 i_2_34 (.ZN (n_96), .A (n_2_2));
NAND2_X1 i_2_33 (.ZN (n_2_1), .A1 (out[32]), .A2 (n_2_36));
AOI222_X1 i_2_32 (.ZN (n_2_0), .A1 (in2[31]), .A2 (CLOCK_slh_n74), .B1 (drc_ipo_n5)
    , .B2 (n_32), .C1 (n_0), .C2 (drc_ipo_n6));
NAND2_X1 i_2_31 (.ZN (n_95), .A1 (n_2_0), .A2 (n_2_1));
MUX2_X1 i_2_30 (.Z (n_94), .A (out[31]), .B (in2[30]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_29 (.Z (n_93), .A (out[30]), .B (in2[29]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_28 (.Z (n_92), .A (out[29]), .B (in2[28]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_27 (.Z (n_91), .A (out[28]), .B (in2[27]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_26 (.Z (n_90), .A (out[27]), .B (in2[26]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_25 (.Z (n_89), .A (out[26]), .B (in2[25]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_24 (.Z (n_88), .A (out[25]), .B (in2[24]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_23 (.Z (n_87), .A (out[24]), .B (in2[23]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_22 (.Z (n_86), .A (out[23]), .B (in2[22]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_21 (.Z (n_85), .A (out[22]), .B (in2[21]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_20 (.Z (n_84), .A (out[21]), .B (in2[20]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_19 (.Z (n_83), .A (out[20]), .B (in2[19]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_18 (.Z (n_82), .A (out[19]), .B (in2[18]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_17 (.Z (n_81), .A (out[18]), .B (in2[17]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_16 (.Z (n_80), .A (out[17]), .B (in2[16]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_15 (.Z (n_79), .A (out[16]), .B (in2[15]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_14 (.Z (n_78), .A (out[15]), .B (in2[14]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_13 (.Z (n_77), .A (out[14]), .B (in2[13]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_12 (.Z (n_76), .A (out[13]), .B (in2[12]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_11 (.Z (n_75), .A (out[12]), .B (in2[11]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_10 (.Z (n_74), .A (out[11]), .B (in2[10]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_9 (.Z (n_73), .A (out[10]), .B (in2[9]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_8 (.Z (n_72), .A (out[9]), .B (in2[8]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_7 (.Z (n_71), .A (out[8]), .B (in2[7]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_6 (.Z (n_70), .A (out[7]), .B (in2[6]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_5 (.Z (n_69), .A (out[6]), .B (in2[5]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_4 (.Z (n_68), .A (out[5]), .B (in2[4]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_3 (.Z (n_67), .A (out[4]), .B (in2[3]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_2 (.Z (n_66), .A (out[3]), .B (in2[2]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_1 (.Z (n_65), .A (out[2]), .B (in2[1]), .S (CLOCK_slh_n74));
MUX2_X1 i_2_0 (.Z (n_64), .A (out[1]), .B (in2[0]), .S (CLOCK_slh_n74));
datapath__0_31 i_1 (.p_0 ({n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
    n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32}), .a ({out[63], uc_1, 
    out[61], out[60], out[59], out[58], out[57], out[56], out[55], out[54], out[53], 
    out[52], out[51], out[50], out[49], out[48], out[47], out[46], out[45], out[44], 
    out[43], out[42], out[41], out[40], out[39], out[38], out[37], out[36], out[35], 
    out[34], out[33], out[32]}), .m ({\m[31] , \m[30] , \m[29] , \m[28] , \m[27] , 
    \m[26] , \m[25] , \m[24] , \m[23] , \m[22] , \m[21] , \m[20] , \m[19] , \m[18] , 
    \m[17] , \m[16] , \m[15] , \m[14] , \m[13] , \m[12] , \m[11] , \m[10] , \m[9] , 
    \m[8] , \m[7] , \m[6] , \m[5] , \m[4] , \m[3] , \m[2] , \m[1] , \m[0] }));
datapath i_0 (.p_0 ({n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, 
    n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, 
    n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}), .a ({out[63], uc_0, out[61], out[60], 
    out[59], out[58], out[57], out[56], out[55], out[54], out[53], out[52], out[51], 
    out[50], out[49], out[48], out[47], out[46], out[45], out[44], out[43], out[42], 
    out[41], out[40], out[39], out[38], out[37], out[36], out[35], out[34], out[33], 
    out[32]}), .m ({\m[31] , \m[30] , \m[29] , \m[28] , \m[27] , \m[26] , \m[25] , 
    \m[24] , \m[23] , \m[22] , \m[21] , \m[20] , \m[19] , \m[18] , \m[17] , \m[16] , 
    \m[15] , \m[14] , \m[13] , \m[12] , \m[11] , \m[10] , \m[9] , \m[8] , \m[7] , 
    \m[6] , \m[5] , \m[4] , \m[3] , \m[2] , \m[1] , \m[0] }));
BUF_X2 drc_ipo_c6 (.Z (drc_ipo_n6), .A (n_2_33));
BUF_X2 drc_ipo_c5 (.Z (drc_ipo_n5), .A (n_2_34));
INV_X4 CTS_L6_c_tid1_13 (.ZN (CTS_n_tid1_14), .A (clk__CTS_1_PP_0));
INV_X4 CTS_L5_c_tid1_24 (.ZN (clk__CTS_1_PP_0), .A (CTS_n_tid1_26));
CLKBUF_X3 CTS_L4_c_tid1_26 (.Z (CTS_n_tid1_26), .A (CTS_n_tid1_29));
INV_X4 CTS_L3_c_tid1_35 (.ZN (CTS_n_tid1_29), .A (CTS_n_tid1_30));
INV_X4 CTS_L2_c_tid1_36 (.ZN (CTS_n_tid1_30), .A (clk__CTS_1_PP_1));
BUF_X16 CLOCK_slh__c50 (.Z (CLOCK_slh_n74), .A (rst));

endmodule //booth_multiplier

module registerNbits (clk__CTS_1_PP_2, clk__CTS_1_PP_27, clk__CTS_1_PP_31, clk, inp, 
    out);

output [31:0] out;
output clk__CTS_1_PP_2;
input clk;
input [31:0] inp;
input clk__CTS_1_PP_27;
input clk__CTS_1_PP_31;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk__CTS_1_PP_2), .D (inp[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk__CTS_1_PP_2), .D (inp[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk__CTS_1_PP_2), .D (inp[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk__CTS_1_PP_2), .D (inp[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk__CTS_1_PP_2), .D (inp[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk__CTS_1_PP_2), .D (inp[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk__CTS_1_PP_2), .D (inp[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk__CTS_1_PP_2), .D (inp[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk__CTS_1_PP_2), .D (inp[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk__CTS_1_PP_2), .D (inp[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk__CTS_1_PP_2), .D (inp[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk__CTS_1_PP_2), .D (inp[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk__CTS_1_PP_2), .D (inp[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk__CTS_1_PP_2), .D (inp[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk__CTS_1_PP_2), .D (inp[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk__CTS_1_PP_27), .D (inp[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk__CTS_1_PP_2), .D (inp[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk__CTS_1_PP_27), .D (inp[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk__CTS_1_PP_27), .D (inp[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk__CTS_1_PP_27), .D (inp[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk__CTS_1_PP_27), .D (inp[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk__CTS_1_PP_27), .D (inp[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk__CTS_1_PP_27), .D (inp[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk__CTS_1_PP_27), .D (inp[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk__CTS_1_PP_27), .D (inp[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk__CTS_1_PP_27), .D (inp[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk__CTS_1_PP_27), .D (inp[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk__CTS_1_PP_27), .D (inp[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk__CTS_1_PP_27), .D (inp[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk__CTS_1_PP_27), .D (inp[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk__CTS_1_PP_27), .D (inp[30]));
INV_X4 CTS_L9_c_tid1_4 (.ZN (clk__CTS_1_PP_2), .A (clk__CTS_1_PP_31));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk__CTS_1_PP_27), .D (inp[31]));

endmodule //registerNbits

module registerNbits__0_102 (clk__CTS_1_PP_2, clk__CTS_1_PP_36, clk__CTS_1_PP_31, 
    clk__CTS_1_PP_37, clk, inp, out);

output [31:0] out;
output clk__CTS_1_PP_2;
output clk__CTS_1_PP_36;
input clk;
input [31:0] inp;
input clk__CTS_1_PP_31;
input clk__CTS_1_PP_37;
wire CTS_n_tid1_184;
wire CTS_n_tid1_186;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk__CTS_1_PP_2), .D (inp[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk__CTS_1_PP_31), .D (inp[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk__CTS_1_PP_31), .D (inp[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk__CTS_1_PP_31), .D (inp[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk__CTS_1_PP_31), .D (inp[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk__CTS_1_PP_31), .D (inp[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk__CTS_1_PP_31), .D (inp[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk__CTS_1_PP_31), .D (inp[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk__CTS_1_PP_31), .D (inp[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk__CTS_1_PP_31), .D (inp[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk__CTS_1_PP_31), .D (inp[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk__CTS_1_PP_31), .D (inp[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk__CTS_1_PP_31), .D (inp[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk__CTS_1_PP_31), .D (inp[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk__CTS_1_PP_31), .D (inp[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk__CTS_1_PP_31), .D (inp[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk__CTS_1_PP_31), .D (inp[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk__CTS_1_PP_2), .D (inp[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk__CTS_1_PP_2), .D (inp[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk__CTS_1_PP_2), .D (inp[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk__CTS_1_PP_2), .D (inp[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk__CTS_1_PP_2), .D (inp[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk__CTS_1_PP_2), .D (inp[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk__CTS_1_PP_2), .D (inp[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk__CTS_1_PP_2), .D (inp[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk__CTS_1_PP_2), .D (inp[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk__CTS_1_PP_2), .D (inp[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk__CTS_1_PP_2), .D (inp[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk__CTS_1_PP_2), .D (inp[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk__CTS_1_PP_2), .D (inp[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk__CTS_1_PP_2), .D (inp[30]));
INV_X16 CTS_L7_c_tid1_23 (.ZN (CTS_n_tid1_184), .A (CTS_n_tid1_186));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk__CTS_1_PP_2), .D (inp[31]));
INV_X4 CTS_L9_c_tid1_6 (.ZN (clk__CTS_1_PP_2), .A (clk__CTS_1_PP_36));
INV_X4 CTS_L8_c_tid1_22 (.ZN (clk__CTS_1_PP_36), .A (CTS_n_tid1_184));
INV_X32 CTS_L6_c_tid1_28 (.ZN (CTS_n_tid1_186), .A (clk__CTS_1_PP_37));

endmodule //registerNbits__0_102

module integrationMult (clk, reset, inputA, inputB, result);

output [63:0] result;
input clk;
input [31:0] inputA;
input [31:0] inputB;
input reset;
wire n_tid1_212;
wire uc_0;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire \outA_reg[63] ;
wire \outA_reg[61] ;
wire \outA_reg[60] ;
wire \outA_reg[59] ;
wire \outA_reg[58] ;
wire \outA_reg[57] ;
wire \outA_reg[56] ;
wire \outA_reg[55] ;
wire \outA_reg[54] ;
wire \outA_reg[53] ;
wire \outA_reg[52] ;
wire \outA_reg[51] ;
wire \outA_reg[50] ;
wire \outA_reg[49] ;
wire \outA_reg[48] ;
wire \outA_reg[47] ;
wire \outA_reg[46] ;
wire \outA_reg[45] ;
wire \outA_reg[44] ;
wire \outA_reg[43] ;
wire \outA_reg[42] ;
wire \outA_reg[41] ;
wire \outA_reg[40] ;
wire \outA_reg[39] ;
wire \outA_reg[38] ;
wire \outA_reg[37] ;
wire \outA_reg[36] ;
wire \outA_reg[35] ;
wire \outA_reg[34] ;
wire \outA_reg[33] ;
wire \outA_reg[32] ;
wire \outA_reg[31] ;
wire \outA_reg[30] ;
wire \outA_reg[29] ;
wire \outA_reg[28] ;
wire \outA_reg[27] ;
wire \outA_reg[26] ;
wire \outA_reg[25] ;
wire \outA_reg[24] ;
wire \outA_reg[23] ;
wire \outA_reg[22] ;
wire \outA_reg[21] ;
wire \outA_reg[20] ;
wire \outA_reg[19] ;
wire \outA_reg[18] ;
wire \outA_reg[17] ;
wire \outA_reg[16] ;
wire \outA_reg[15] ;
wire \outA_reg[14] ;
wire \outA_reg[13] ;
wire \outA_reg[12] ;
wire \outA_reg[11] ;
wire \outA_reg[10] ;
wire \outA_reg[9] ;
wire \outA_reg[8] ;
wire \outA_reg[7] ;
wire \outA_reg[6] ;
wire \outA_reg[5] ;
wire \outA_reg[4] ;
wire \outA_reg[3] ;
wire \outA_reg[2] ;
wire \outA_reg[1] ;
wire \outA_reg[0] ;
wire uc_1;
wire uc_2;
wire CTS_n_tid1_130;
wire CTS_n_tid1_11;
wire CTS_n_tid1_12;
wire CTS_n_tid1_129;
wire CTS_n_tid1_108;
wire CTS_n_tid1_109;

// WARNING . Detected multiport output net(s). Introducing ASSIGN statements.
// This may cause simulation/synthesis mismatches . 
assign result[63] = result[62];

registerNbits__parameterized0 outB (.out ({result[62], uc_2, result[61], result[60], 
    result[59], result[58], result[57], result[56], result[55], result[54], result[53], 
    result[52], result[51], result[50], result[49], result[48], result[47], result[46], 
    result[45], result[44], result[43], result[42], result[41], result[40], result[39], 
    result[38], result[37], result[36], result[35], result[34], result[33], result[32], 
    result[31], result[30], result[29], result[28], result[27], result[26], result[25], 
    result[24], result[23], result[22], result[21], result[20], result[19], result[18], 
    result[17], result[16], result[15], result[14], result[13], result[12], result[11], 
    result[10], result[9], result[8], result[7], result[6], result[5], result[4], 
    result[3], result[2], result[1], result[0]}), .clk__CTS_1_PP_35 (CTS_n_tid1_108)
    , .clk__CTS_1_PP_36 (CTS_n_tid1_109), .inp ({\outA_reg[63] , uc_1, \outA_reg[61] , 
    \outA_reg[60] , \outA_reg[59] , \outA_reg[58] , \outA_reg[57] , \outA_reg[56] , 
    \outA_reg[55] , \outA_reg[54] , \outA_reg[53] , \outA_reg[52] , \outA_reg[51] , 
    \outA_reg[50] , \outA_reg[49] , \outA_reg[48] , \outA_reg[47] , \outA_reg[46] , 
    \outA_reg[45] , \outA_reg[44] , \outA_reg[43] , \outA_reg[42] , \outA_reg[41] , 
    \outA_reg[40] , \outA_reg[39] , \outA_reg[38] , \outA_reg[37] , \outA_reg[36] , 
    \outA_reg[35] , \outA_reg[34] , \outA_reg[33] , \outA_reg[32] , \outA_reg[31] , 
    \outA_reg[30] , \outA_reg[29] , \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , 
    \outA_reg[25] , \outA_reg[24] , \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , 
    \outA_reg[20] , \outA_reg[19] , \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , 
    \outA_reg[15] , \outA_reg[14] , \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , 
    \outA_reg[10] , \outA_reg[9] , \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , 
    \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , \outA_reg[1] , \outA_reg[0] }), .clk__CTS_1_PP_2 (CTS_n_tid1_11)
    , .clk__CTS_1_PP_3 (CTS_n_tid1_12), .clk__CTS_1_PP_41 (CTS_n_tid1_129));
booth_multiplier mult (.out ({\outA_reg[63] , uc_0, \outA_reg[61] , \outA_reg[60] , 
    \outA_reg[59] , \outA_reg[58] , \outA_reg[57] , \outA_reg[56] , \outA_reg[55] , 
    \outA_reg[54] , \outA_reg[53] , \outA_reg[52] , \outA_reg[51] , \outA_reg[50] , 
    \outA_reg[49] , \outA_reg[48] , \outA_reg[47] , \outA_reg[46] , \outA_reg[45] , 
    \outA_reg[44] , \outA_reg[43] , \outA_reg[42] , \outA_reg[41] , \outA_reg[40] , 
    \outA_reg[39] , \outA_reg[38] , \outA_reg[37] , \outA_reg[36] , \outA_reg[35] , 
    \outA_reg[34] , \outA_reg[33] , \outA_reg[32] , \outA_reg[31] , \outA_reg[30] , 
    \outA_reg[29] , \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , 
    \outA_reg[24] , \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , 
    \outA_reg[19] , \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , 
    \outA_reg[14] , \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , 
    \outA_reg[9] , \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , 
    \outA_reg[3] , \outA_reg[2] , \outA_reg[1] , \outA_reg[0] }), .clk__CTS_1_PP_0 (CTS_n_tid1_130)
    , .in1 ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , \A_reg[27] , \A_reg[26] , 
    \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , \A_reg[21] , \A_reg[20] , 
    \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , \A_reg[15] , \A_reg[14] , 
    \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , \A_reg[9] , \A_reg[8] , \A_reg[7] , 
    \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , \A_reg[1] , \A_reg[0] })
    , .in2 ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , \B_reg[26] , 
    \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , \B_reg[20] , 
    \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , \B_reg[14] , 
    \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , \B_reg[8] , \B_reg[7] , 
    \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] })
    , .rst (reset), .clk__CTS_1_PP_1 (n_tid1_212));
registerNbits regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , 
    \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , 
    \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , 
    \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , 
    \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , 
    \B_reg[1] , \B_reg[0] }), .clk__CTS_1_PP_2 (CTS_n_tid1_12), .inp ({inputB[31], 
    inputB[30], inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], inputB[24], 
    inputB[23], inputB[22], inputB[21], inputB[20], inputB[19], inputB[18], inputB[17], 
    inputB[16], inputB[15], inputB[14], inputB[13], inputB[12], inputB[11], inputB[10], 
    inputB[9], inputB[8], inputB[7], inputB[6], inputB[5], inputB[4], inputB[3], 
    inputB[2], inputB[1], inputB[0]}), .clk__CTS_1_PP_27 (CTS_n_tid1_109), .clk__CTS_1_PP_31 (CTS_n_tid1_129));
registerNbits__0_102 regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .clk__CTS_1_PP_2 (CTS_n_tid1_11), .clk__CTS_1_PP_36 (CTS_n_tid1_129)
    , .inp ({inputA[31], inputA[30], inputA[29], inputA[28], inputA[27], inputA[26], 
    inputA[25], inputA[24], inputA[23], inputA[22], inputA[21], inputA[20], inputA[19], 
    inputA[18], inputA[17], inputA[16], inputA[15], inputA[14], inputA[13], inputA[12], 
    inputA[11], inputA[10], inputA[9], inputA[8], inputA[7], inputA[6], inputA[5], 
    inputA[4], inputA[3], inputA[2], inputA[1], inputA[0]}), .clk__CTS_1_PP_31 (CTS_n_tid1_108), .clk__CTS_1_PP_37 (CTS_n_tid1_130));
BUF_X8 CTS_L1_tid1__c1_tid1__c57 (.Z (n_tid1_212), .A (clk));

endmodule //integrationMult


