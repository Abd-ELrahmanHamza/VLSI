/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 23 14:35:33 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2003289718 */

module registerNbits__0_22(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits__0_25(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module datapath(p_0, in2);
   output [31:0]p_0;
   input [31:0]in2;

   XOR2_X1 i_0 (.A(in2[1]), .B(in2[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(in2[2]), .B1(in2[1]), .B2(in2[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(in2[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(in2[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(in2[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(in2[6]), .B1(n_27), .B2(in2[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(in2[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(in2[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(in2[9]), .B1(n_25), .B2(in2[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(in2[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(in2[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(in2[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(in2[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(in2[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(in2[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(in2[16]), .B1(n_19), .B2(in2[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(in2[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(in2[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(in2[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(in2[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(in2[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(in2[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(in2[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(in2[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(in2[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(in2[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(in2[27]), .B1(n_9), .B2(in2[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(in2[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(in2[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(in2[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(in2[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(in2[28]), .A3(in2[29]), .A4(in2[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(in2[28]), .A3(in2[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(in2[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(in2[26]), .A3(in2[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(in2[23]), .A3(in2[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(in2[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(in2[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(in2[18]), .A3(in2[19]), .A4(in2[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(in2[18]), .A3(in2[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(in2[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(in2[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(in2[15]), .A3(in2[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(in2[12]), .A3(in2[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(in2[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(in2[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(in2[8]), .A3(in2[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(in2[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(in2[5]), .A3(in2[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(in2[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(in2[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(in2[2]), .A2(in2[1]), .A3(in2[0]), .ZN(n_29));
   INV_X1 i_61 (.A(in2[11]), .ZN(n_30));
   INV_X1 i_62 (.A(in2[14]), .ZN(n_31));
   INV_X1 i_63 (.A(in2[21]), .ZN(n_32));
   INV_X1 i_64 (.A(in2[25]), .ZN(n_33));
endmodule

module datapath__0_2(p_0, in1);
   output [31:0]p_0;
   input [31:0]in1;

   XOR2_X1 i_0 (.A(in1[1]), .B(in1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(in1[2]), .B1(in1[1]), .B2(in1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(in1[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(in1[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(in1[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(in1[6]), .B1(n_27), .B2(in1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(in1[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(in1[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(in1[9]), .B1(n_25), .B2(in1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(in1[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(in1[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(in1[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(in1[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(in1[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(in1[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(in1[16]), .B1(n_19), .B2(in1[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(in1[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(in1[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(in1[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(in1[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(in1[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(in1[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(in1[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(in1[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(in1[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(in1[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(in1[27]), .B1(n_9), .B2(in1[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(in1[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(in1[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(in1[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(in1[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(in1[28]), .A3(in1[29]), .A4(in1[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(in1[28]), .A3(in1[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(in1[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(in1[26]), .A3(in1[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(in1[23]), .A3(in1[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(in1[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(in1[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(in1[18]), .A3(in1[19]), .A4(in1[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(in1[18]), .A3(in1[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(in1[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(in1[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(in1[15]), .A3(in1[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(in1[12]), .A3(in1[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(in1[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(in1[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(in1[8]), .A3(in1[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(in1[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(in1[5]), .A3(in1[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(in1[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(in1[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(in1[2]), .A2(in1[1]), .A3(in1[0]), .ZN(n_29));
   INV_X1 i_61 (.A(in1[11]), .ZN(n_30));
   INV_X1 i_62 (.A(in1[14]), .ZN(n_31));
   INV_X1 i_63 (.A(in1[21]), .ZN(n_32));
   INV_X1 i_64 (.A(in1[25]), .ZN(n_33));
endmodule

module datapath__0_9(m, p_0, p_1);
   input [31:0]m;
   input [31:0]p_0;
   output [32:0]p_1;

   HA_X1 i_0 (.A(m[0]), .B(p_0[0]), .CO(n_0), .S(p_1[0]));
   FA_X1 i_1 (.A(m[1]), .B(p_0[1]), .CI(n_0), .CO(n_1), .S(p_1[1]));
   FA_X1 i_2 (.A(m[2]), .B(p_0[2]), .CI(n_1), .CO(n_2), .S(p_1[2]));
   FA_X1 i_3 (.A(m[3]), .B(p_0[3]), .CI(n_2), .CO(n_3), .S(p_1[3]));
   FA_X1 i_4 (.A(m[4]), .B(p_0[4]), .CI(n_3), .CO(n_4), .S(p_1[4]));
   FA_X1 i_5 (.A(m[5]), .B(p_0[5]), .CI(n_4), .CO(n_5), .S(p_1[5]));
   FA_X1 i_6 (.A(m[6]), .B(p_0[6]), .CI(n_5), .CO(n_6), .S(p_1[6]));
   FA_X1 i_7 (.A(m[7]), .B(p_0[7]), .CI(n_6), .CO(n_7), .S(p_1[7]));
   FA_X1 i_8 (.A(m[8]), .B(p_0[8]), .CI(n_7), .CO(n_8), .S(p_1[8]));
   FA_X1 i_9 (.A(m[9]), .B(p_0[9]), .CI(n_8), .CO(n_9), .S(p_1[9]));
   FA_X1 i_10 (.A(m[10]), .B(p_0[10]), .CI(n_9), .CO(n_10), .S(p_1[10]));
   FA_X1 i_11 (.A(m[11]), .B(p_0[11]), .CI(n_10), .CO(n_11), .S(p_1[11]));
   FA_X1 i_12 (.A(m[12]), .B(p_0[12]), .CI(n_11), .CO(n_12), .S(p_1[12]));
   FA_X1 i_13 (.A(m[13]), .B(p_0[13]), .CI(n_12), .CO(n_13), .S(p_1[13]));
   FA_X1 i_14 (.A(m[14]), .B(p_0[14]), .CI(n_13), .CO(n_14), .S(p_1[14]));
   FA_X1 i_15 (.A(m[15]), .B(p_0[15]), .CI(n_14), .CO(n_15), .S(p_1[15]));
   FA_X1 i_16 (.A(m[16]), .B(p_0[16]), .CI(n_15), .CO(n_16), .S(p_1[16]));
   FA_X1 i_17 (.A(m[17]), .B(p_0[17]), .CI(n_16), .CO(n_17), .S(p_1[17]));
   FA_X1 i_18 (.A(m[18]), .B(p_0[18]), .CI(n_17), .CO(n_18), .S(p_1[18]));
   FA_X1 i_19 (.A(m[19]), .B(p_0[19]), .CI(n_18), .CO(n_19), .S(p_1[19]));
   FA_X1 i_20 (.A(m[20]), .B(p_0[20]), .CI(n_19), .CO(n_20), .S(p_1[20]));
   FA_X1 i_21 (.A(m[21]), .B(p_0[21]), .CI(n_20), .CO(n_21), .S(p_1[21]));
   FA_X1 i_22 (.A(m[22]), .B(p_0[22]), .CI(n_21), .CO(n_22), .S(p_1[22]));
   FA_X1 i_23 (.A(m[23]), .B(p_0[23]), .CI(n_22), .CO(n_23), .S(p_1[23]));
   FA_X1 i_24 (.A(m[24]), .B(p_0[24]), .CI(n_23), .CO(n_24), .S(p_1[24]));
   FA_X1 i_25 (.A(m[25]), .B(p_0[25]), .CI(n_24), .CO(n_25), .S(p_1[25]));
   FA_X1 i_26 (.A(m[26]), .B(p_0[26]), .CI(n_25), .CO(n_26), .S(p_1[26]));
   FA_X1 i_27 (.A(m[27]), .B(p_0[27]), .CI(n_26), .CO(n_27), .S(p_1[27]));
   FA_X1 i_28 (.A(m[28]), .B(p_0[28]), .CI(n_27), .CO(n_28), .S(p_1[28]));
   FA_X1 i_29 (.A(m[29]), .B(p_0[29]), .CI(n_28), .CO(n_29), .S(p_1[29]));
   FA_X1 i_30 (.A(m[30]), .B(p_0[30]), .CI(n_29), .CO(n_30), .S(p_1[30]));
   FA_X1 i_31 (.A(m[31]), .B(p_0[31]), .CI(n_30), .CO(p_1[32]), .S(p_1[31]));
endmodule

module datapath__0_11(p_0, p_1);
   output [64:0]p_0;
   input [64:0]p_1;

   XOR2_X1 i_0 (.A(p_1[1]), .B(p_1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_61), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(p_1[2]), .B1(p_1[1]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[3]), .B(n_61), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(p_1[4]), .B(n_60), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(p_1[5]), .B(n_59), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_58), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(p_1[6]), .B1(n_59), .B2(p_1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[7]), .B(n_58), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(p_1[8]), .B(n_57), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_56), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(p_1[9]), .B1(n_57), .B2(p_1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[10]), .B(n_56), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(p_1[11]), .B(n_55), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(p_1[12]), .B(n_54), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(p_1[13]), .B(n_53), .ZN(p_0[13]));
   XOR2_X1 i_16 (.A(p_1[14]), .B(n_52), .Z(p_0[14]));
   AND2_X1 i_17 (.A1(n_51), .A2(n_3), .ZN(p_0[15]));
   OAI21_X1 i_18 (.A(p_1[15]), .B1(n_52), .B2(p_1[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(p_1[16]), .B(n_51), .Z(p_0[16]));
   XOR2_X1 i_20 (.A(p_1[17]), .B(n_50), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(p_1[18]), .B(n_49), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(p_1[19]), .B(n_48), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(p_1[20]), .B(n_47), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(p_1[21]), .B(n_46), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(p_1[22]), .B(n_45), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(p_1[23]), .B(n_44), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(p_1[24]), .B(n_43), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(p_1[25]), .B(n_42), .ZN(p_0[25]));
   XNOR2_X1 i_29 (.A(p_1[26]), .B(n_41), .ZN(p_0[26]));
   XOR2_X1 i_30 (.A(p_1[27]), .B(n_40), .Z(p_0[27]));
   XOR2_X1 i_31 (.A(p_1[28]), .B(n_39), .Z(p_0[28]));
   XNOR2_X1 i_32 (.A(p_1[29]), .B(n_38), .ZN(p_0[29]));
   XNOR2_X1 i_33 (.A(p_1[30]), .B(n_37), .ZN(p_0[30]));
   XNOR2_X1 i_34 (.A(p_1[31]), .B(n_36), .ZN(p_0[31]));
   XOR2_X1 i_35 (.A(p_1[32]), .B(n_35), .Z(p_0[32]));
   XOR2_X1 i_36 (.A(p_1[33]), .B(n_34), .Z(p_0[33]));
   XNOR2_X1 i_37 (.A(p_1[34]), .B(n_33), .ZN(p_0[34]));
   XNOR2_X1 i_38 (.A(p_1[35]), .B(n_32), .ZN(p_0[35]));
   XNOR2_X1 i_39 (.A(p_1[36]), .B(n_31), .ZN(p_0[36]));
   XOR2_X1 i_40 (.A(p_1[37]), .B(n_30), .Z(p_0[37]));
   XOR2_X1 i_41 (.A(p_1[38]), .B(n_29), .Z(p_0[38]));
   XNOR2_X1 i_42 (.A(p_1[39]), .B(n_28), .ZN(p_0[39]));
   XNOR2_X1 i_43 (.A(p_1[40]), .B(n_27), .ZN(p_0[40]));
   XOR2_X1 i_44 (.A(p_1[41]), .B(n_26), .Z(p_0[41]));
   XNOR2_X1 i_45 (.A(p_1[42]), .B(n_25), .ZN(p_0[42]));
   XOR2_X1 i_46 (.A(p_1[43]), .B(n_24), .Z(p_0[43]));
   AND2_X1 i_47 (.A1(n_23), .A2(n_4), .ZN(p_0[44]));
   OAI21_X1 i_48 (.A(p_1[44]), .B1(n_24), .B2(p_1[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(p_1[45]), .B(n_23), .Z(p_0[45]));
   XOR2_X1 i_50 (.A(p_1[46]), .B(n_22), .Z(p_0[46]));
   XOR2_X1 i_51 (.A(p_1[47]), .B(n_21), .Z(p_0[47]));
   XOR2_X1 i_52 (.A(p_1[48]), .B(n_20), .Z(p_0[48]));
   XNOR2_X1 i_53 (.A(p_1[49]), .B(n_19), .ZN(p_0[49]));
   XNOR2_X1 i_54 (.A(p_1[50]), .B(n_18), .ZN(p_0[50]));
   XNOR2_X1 i_55 (.A(p_1[51]), .B(n_17), .ZN(p_0[51]));
   XOR2_X1 i_56 (.A(p_1[52]), .B(n_16), .Z(p_0[52]));
   XNOR2_X1 i_57 (.A(p_1[53]), .B(n_15), .ZN(p_0[53]));
   XNOR2_X1 i_58 (.A(p_1[54]), .B(n_14), .ZN(p_0[54]));
   XNOR2_X1 i_59 (.A(p_1[55]), .B(n_13), .ZN(p_0[55]));
   XOR2_X1 i_60 (.A(p_1[56]), .B(n_12), .Z(p_0[56]));
   AND2_X1 i_61 (.A1(n_11), .A2(n_5), .ZN(p_0[57]));
   OAI21_X1 i_62 (.A(p_1[57]), .B1(n_12), .B2(p_1[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(p_1[58]), .B(n_11), .Z(p_0[58]));
   XNOR2_X1 i_64 (.A(p_1[59]), .B(n_10), .ZN(p_0[59]));
   XNOR2_X1 i_65 (.A(p_1[60]), .B(n_9), .ZN(p_0[60]));
   XOR2_X1 i_66 (.A(p_1[61]), .B(n_8), .Z(p_0[61]));
   XNOR2_X1 i_67 (.A(p_1[62]), .B(n_7), .ZN(p_0[62]));
   XNOR2_X1 i_68 (.A(p_1[63]), .B(n_6), .ZN(p_0[63]));
   NAND2_X1 i_69 (.A1(n_6), .A2(n_73), .ZN(p_0[64]));
   NOR3_X1 i_70 (.A1(n_8), .A2(p_1[61]), .A3(p_1[62]), .ZN(n_6));
   NOR2_X1 i_71 (.A1(n_8), .A2(p_1[61]), .ZN(n_7));
   NAND2_X1 i_72 (.A1(n_9), .A2(n_72), .ZN(n_8));
   NOR3_X1 i_73 (.A1(n_11), .A2(p_1[58]), .A3(p_1[59]), .ZN(n_9));
   NOR2_X1 i_74 (.A1(n_11), .A2(p_1[58]), .ZN(n_10));
   OR3_X1 i_75 (.A1(n_12), .A2(p_1[56]), .A3(p_1[57]), .ZN(n_11));
   NAND2_X1 i_76 (.A1(n_13), .A2(n_71), .ZN(n_12));
   NOR4_X1 i_77 (.A1(n_16), .A2(p_1[52]), .A3(p_1[53]), .A4(p_1[54]), .ZN(n_13));
   NOR3_X1 i_78 (.A1(n_16), .A2(p_1[52]), .A3(p_1[53]), .ZN(n_14));
   NOR2_X1 i_79 (.A1(n_16), .A2(p_1[52]), .ZN(n_15));
   NAND2_X1 i_80 (.A1(n_17), .A2(n_70), .ZN(n_16));
   NOR4_X1 i_81 (.A1(n_20), .A2(p_1[48]), .A3(p_1[49]), .A4(p_1[50]), .ZN(n_17));
   NOR3_X1 i_82 (.A1(n_20), .A2(p_1[48]), .A3(p_1[49]), .ZN(n_18));
   NOR2_X1 i_83 (.A1(n_20), .A2(p_1[48]), .ZN(n_19));
   OR2_X1 i_84 (.A1(n_21), .A2(p_1[47]), .ZN(n_20));
   OR2_X1 i_85 (.A1(n_22), .A2(p_1[46]), .ZN(n_21));
   OR2_X1 i_86 (.A1(n_23), .A2(p_1[45]), .ZN(n_22));
   OR3_X1 i_87 (.A1(n_24), .A2(p_1[43]), .A3(p_1[44]), .ZN(n_23));
   NAND2_X1 i_88 (.A1(n_25), .A2(n_69), .ZN(n_24));
   NOR2_X1 i_89 (.A1(n_26), .A2(p_1[41]), .ZN(n_25));
   NAND2_X1 i_90 (.A1(n_27), .A2(n_68), .ZN(n_26));
   NOR3_X1 i_91 (.A1(n_29), .A2(p_1[38]), .A3(p_1[39]), .ZN(n_27));
   NOR2_X1 i_92 (.A1(n_29), .A2(p_1[38]), .ZN(n_28));
   OR2_X1 i_93 (.A1(n_30), .A2(p_1[37]), .ZN(n_29));
   NAND2_X1 i_94 (.A1(n_31), .A2(n_67), .ZN(n_30));
   NOR4_X1 i_95 (.A1(n_34), .A2(p_1[33]), .A3(p_1[34]), .A4(p_1[35]), .ZN(n_31));
   NOR3_X1 i_96 (.A1(n_34), .A2(p_1[33]), .A3(p_1[34]), .ZN(n_32));
   NOR2_X1 i_97 (.A1(n_34), .A2(p_1[33]), .ZN(n_33));
   OR2_X1 i_98 (.A1(n_35), .A2(p_1[32]), .ZN(n_34));
   NAND2_X1 i_99 (.A1(n_36), .A2(n_66), .ZN(n_35));
   NOR4_X1 i_100 (.A1(n_39), .A2(p_1[28]), .A3(p_1[29]), .A4(p_1[30]), .ZN(n_36));
   NOR3_X1 i_101 (.A1(n_39), .A2(p_1[28]), .A3(p_1[29]), .ZN(n_37));
   NOR2_X1 i_102 (.A1(n_39), .A2(p_1[28]), .ZN(n_38));
   OR2_X1 i_103 (.A1(n_40), .A2(p_1[27]), .ZN(n_39));
   NAND2_X1 i_104 (.A1(n_41), .A2(n_65), .ZN(n_40));
   NOR4_X1 i_105 (.A1(n_44), .A2(p_1[23]), .A3(p_1[24]), .A4(p_1[25]), .ZN(n_41));
   NOR3_X1 i_106 (.A1(n_44), .A2(p_1[23]), .A3(p_1[24]), .ZN(n_42));
   NOR2_X1 i_107 (.A1(n_44), .A2(p_1[23]), .ZN(n_43));
   OR2_X1 i_108 (.A1(n_45), .A2(p_1[22]), .ZN(n_44));
   NAND2_X1 i_109 (.A1(n_46), .A2(n_64), .ZN(n_45));
   NOR4_X1 i_110 (.A1(n_49), .A2(p_1[18]), .A3(p_1[19]), .A4(p_1[20]), .ZN(n_46));
   NOR3_X1 i_111 (.A1(n_49), .A2(p_1[18]), .A3(p_1[19]), .ZN(n_47));
   NOR2_X1 i_112 (.A1(n_49), .A2(p_1[18]), .ZN(n_48));
   OR2_X1 i_113 (.A1(n_50), .A2(p_1[17]), .ZN(n_49));
   OR2_X1 i_114 (.A1(n_51), .A2(p_1[16]), .ZN(n_50));
   OR3_X1 i_115 (.A1(n_52), .A2(p_1[14]), .A3(p_1[15]), .ZN(n_51));
   NAND2_X1 i_116 (.A1(n_53), .A2(n_63), .ZN(n_52));
   NOR2_X1 i_117 (.A1(n_54), .A2(p_1[12]), .ZN(n_53));
   NAND2_X1 i_118 (.A1(n_55), .A2(n_62), .ZN(n_54));
   NOR2_X1 i_119 (.A1(n_56), .A2(p_1[10]), .ZN(n_55));
   OR3_X1 i_120 (.A1(n_57), .A2(p_1[8]), .A3(p_1[9]), .ZN(n_56));
   OR2_X1 i_121 (.A1(n_58), .A2(p_1[7]), .ZN(n_57));
   OR3_X1 i_122 (.A1(n_59), .A2(p_1[5]), .A3(p_1[6]), .ZN(n_58));
   OR2_X1 i_123 (.A1(n_60), .A2(p_1[4]), .ZN(n_59));
   OR2_X1 i_124 (.A1(n_61), .A2(p_1[3]), .ZN(n_60));
   OR3_X1 i_125 (.A1(p_1[2]), .A2(p_1[1]), .A3(p_1[0]), .ZN(n_61));
   INV_X1 i_126 (.A(p_1[11]), .ZN(n_62));
   INV_X1 i_127 (.A(p_1[13]), .ZN(n_63));
   INV_X1 i_128 (.A(p_1[21]), .ZN(n_64));
   INV_X1 i_129 (.A(p_1[26]), .ZN(n_65));
   INV_X1 i_130 (.A(p_1[31]), .ZN(n_66));
   INV_X1 i_131 (.A(p_1[36]), .ZN(n_67));
   INV_X1 i_132 (.A(p_1[40]), .ZN(n_68));
   INV_X1 i_133 (.A(p_1[42]), .ZN(n_69));
   INV_X1 i_134 (.A(p_1[51]), .ZN(n_70));
   INV_X1 i_135 (.A(p_1[55]), .ZN(n_71));
   INV_X1 i_136 (.A(p_1[60]), .ZN(n_72));
   INV_X1 i_137 (.A(p_1[63]), .ZN(n_73));
endmodule

module sequentialmultiplier(in1, in2, clk, reset, en, result, enableOutput);
   input [31:0]in1;
   input [31:0]in2;
   input clk;
   input reset;
   input en;
   output [63:0]result;
   output enableOutput;

   wire [5:0]counter;
   wire resetReg;
   wire [64:0]res;
   wire n_1_3;
   wire n_1_0;
   wire n_1_4;
   wire n_1_1;
   wire n_1_5;
   wire n_1_2;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_115;
   wire n_1_116;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_123;
   wire n_1_124;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_149;
   wire n_1_150;
   wire n_1_151;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_160;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_169;
   wire n_1_170;
   wire n_1_171;
   wire n_1_184;
   wire [31:0]m;
   wire n_1_188;
   wire n_1_82;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;
   wire n_1_176;
   wire n_1_177;
   wire n_1_178;
   wire n_1_179;
   wire n_1_180;
   wire n_1_181;
   wire n_1_182;
   wire n_1_183;
   wire n_1_185;
   wire n_1_186;
   wire n_1_187;
   wire n_1_189;

   datapath i_0 (.p_0({n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
      n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, 
      n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, uc_0}), .in2(in2));
   datapath__0_2 i_2 (.p_0({n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, 
      n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, 
      n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, uc_1}), 
      .in1(in1));
   DFF_X1 enableOutput_reg (.D(n_334), .CK(clk), .Q(enableOutput), .QN());
   datapath__0_9 i_9 (.m({m[31], m[30], m[29], m[28], m[27], m[26], m[25], m[24], 
      m[23], m[22], m[21], m[20], m[19], m[18], m[17], m[16], m[15], m[14], 
      m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], 
      m[1], in1[0]}), .p_0({res[63], res[62], res[61], res[60], res[59], res[58], 
      res[57], res[56], res[55], res[54], res[53], res[52], res[51], res[50], 
      res[49], res[48], res[47], res[46], res[45], res[44], res[43], res[42], 
      res[41], res[40], res[39], res[38], res[37], res[36], res[35], res[34], 
      res[33], res[32]}), .p_1({n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
      n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, 
      n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, 
      n_65}));
   datapath__0_11 i_11 (.p_0({n_161, n_160, n_159, n_158, n_157, n_156, n_155, 
      n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, 
      n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, 
      n_134, n_133, n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, 
      n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, 
      n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, 
      n_104, n_103, n_102, n_101, n_100, n_99, n_98, uc_2}), .p_1({1'b0, n_331, 
      n_330, n_329, n_328, n_327, n_326, n_325, n_324, n_323, n_322, n_321, 
      n_320, n_319, n_318, n_317, n_316, n_315, n_314, n_313, n_312, n_311, 
      n_310, n_309, n_308, n_307, n_306, n_305, n_304, n_303, n_302, n_301, 
      n_300, n_299, res[31], res[30], res[29], res[28], res[27], res[26], 
      res[25], res[24], res[23], res[22], res[21], res[20], res[19], res[18], 
      res[17], res[16], res[15], res[14], res[13], res[12], res[11], res[10], 
      res[9], res[8], res[7], res[6], res[5], res[4], res[3], res[2], res[1]}));
   CLKGATETST_X1 clk_gate_result_reg (.CK(clk), .E(n_333), .SE(1'b0), .GCK(n_0));
   DFF_X1 \result_reg[63]  (.D(n_227), .CK(n_0), .Q(result[63]), .QN());
   DFF_X1 \result_reg[62]  (.D(n_226), .CK(n_0), .Q(result[62]), .QN());
   DFF_X1 \result_reg[61]  (.D(n_225), .CK(n_0), .Q(result[61]), .QN());
   DFF_X1 \result_reg[60]  (.D(n_224), .CK(n_0), .Q(result[60]), .QN());
   DFF_X1 \result_reg[59]  (.D(n_223), .CK(n_0), .Q(result[59]), .QN());
   DFF_X1 \result_reg[58]  (.D(n_222), .CK(n_0), .Q(result[58]), .QN());
   DFF_X1 \result_reg[57]  (.D(n_221), .CK(n_0), .Q(result[57]), .QN());
   DFF_X1 \result_reg[56]  (.D(n_220), .CK(n_0), .Q(result[56]), .QN());
   DFF_X1 \result_reg[55]  (.D(n_219), .CK(n_0), .Q(result[55]), .QN());
   DFF_X1 \result_reg[54]  (.D(n_218), .CK(n_0), .Q(result[54]), .QN());
   DFF_X1 \result_reg[53]  (.D(n_217), .CK(n_0), .Q(result[53]), .QN());
   DFF_X1 \result_reg[52]  (.D(n_216), .CK(n_0), .Q(result[52]), .QN());
   DFF_X1 \result_reg[51]  (.D(n_215), .CK(n_0), .Q(result[51]), .QN());
   DFF_X1 \result_reg[50]  (.D(n_214), .CK(n_0), .Q(result[50]), .QN());
   DFF_X1 \result_reg[49]  (.D(n_213), .CK(n_0), .Q(result[49]), .QN());
   DFF_X1 \result_reg[48]  (.D(n_212), .CK(n_0), .Q(result[48]), .QN());
   DFF_X1 \result_reg[47]  (.D(n_211), .CK(n_0), .Q(result[47]), .QN());
   DFF_X1 \result_reg[46]  (.D(n_210), .CK(n_0), .Q(result[46]), .QN());
   DFF_X1 \result_reg[45]  (.D(n_209), .CK(n_0), .Q(result[45]), .QN());
   DFF_X1 \result_reg[44]  (.D(n_208), .CK(n_0), .Q(result[44]), .QN());
   DFF_X1 \result_reg[43]  (.D(n_207), .CK(n_0), .Q(result[43]), .QN());
   DFF_X1 \result_reg[42]  (.D(n_206), .CK(n_0), .Q(result[42]), .QN());
   DFF_X1 \result_reg[41]  (.D(n_205), .CK(n_0), .Q(result[41]), .QN());
   DFF_X1 \result_reg[40]  (.D(n_204), .CK(n_0), .Q(result[40]), .QN());
   DFF_X1 \result_reg[39]  (.D(n_203), .CK(n_0), .Q(result[39]), .QN());
   DFF_X1 \result_reg[38]  (.D(n_202), .CK(n_0), .Q(result[38]), .QN());
   DFF_X1 \result_reg[37]  (.D(n_201), .CK(n_0), .Q(result[37]), .QN());
   DFF_X1 \result_reg[36]  (.D(n_200), .CK(n_0), .Q(result[36]), .QN());
   DFF_X1 \result_reg[35]  (.D(n_199), .CK(n_0), .Q(result[35]), .QN());
   DFF_X1 \result_reg[34]  (.D(n_198), .CK(n_0), .Q(result[34]), .QN());
   DFF_X1 \result_reg[33]  (.D(n_197), .CK(n_0), .Q(result[33]), .QN());
   DFF_X1 \result_reg[32]  (.D(n_196), .CK(n_0), .Q(result[32]), .QN());
   DFF_X1 \result_reg[31]  (.D(n_195), .CK(n_0), .Q(result[31]), .QN());
   DFF_X1 \result_reg[30]  (.D(n_194), .CK(n_0), .Q(result[30]), .QN());
   DFF_X1 \result_reg[29]  (.D(n_193), .CK(n_0), .Q(result[29]), .QN());
   DFF_X1 \result_reg[28]  (.D(n_192), .CK(n_0), .Q(result[28]), .QN());
   DFF_X1 \result_reg[27]  (.D(n_191), .CK(n_0), .Q(result[27]), .QN());
   DFF_X1 \result_reg[26]  (.D(n_190), .CK(n_0), .Q(result[26]), .QN());
   DFF_X1 \result_reg[25]  (.D(n_189), .CK(n_0), .Q(result[25]), .QN());
   DFF_X1 \result_reg[24]  (.D(n_188), .CK(n_0), .Q(result[24]), .QN());
   DFF_X1 \result_reg[23]  (.D(n_187), .CK(n_0), .Q(result[23]), .QN());
   DFF_X1 \result_reg[22]  (.D(n_186), .CK(n_0), .Q(result[22]), .QN());
   DFF_X1 \result_reg[21]  (.D(n_185), .CK(n_0), .Q(result[21]), .QN());
   DFF_X1 \result_reg[20]  (.D(n_184), .CK(n_0), .Q(result[20]), .QN());
   DFF_X1 \result_reg[19]  (.D(n_183), .CK(n_0), .Q(result[19]), .QN());
   DFF_X1 \result_reg[18]  (.D(n_182), .CK(n_0), .Q(result[18]), .QN());
   DFF_X1 \result_reg[17]  (.D(n_181), .CK(n_0), .Q(result[17]), .QN());
   DFF_X1 \result_reg[16]  (.D(n_180), .CK(n_0), .Q(result[16]), .QN());
   DFF_X1 \result_reg[15]  (.D(n_179), .CK(n_0), .Q(result[15]), .QN());
   DFF_X1 \result_reg[14]  (.D(n_178), .CK(n_0), .Q(result[14]), .QN());
   DFF_X1 \result_reg[13]  (.D(n_177), .CK(n_0), .Q(result[13]), .QN());
   DFF_X1 \result_reg[12]  (.D(n_176), .CK(n_0), .Q(result[12]), .QN());
   DFF_X1 \result_reg[11]  (.D(n_175), .CK(n_0), .Q(result[11]), .QN());
   DFF_X1 \result_reg[10]  (.D(n_174), .CK(n_0), .Q(result[10]), .QN());
   DFF_X1 \result_reg[9]  (.D(n_173), .CK(n_0), .Q(result[9]), .QN());
   DFF_X1 \result_reg[8]  (.D(n_172), .CK(n_0), .Q(result[8]), .QN());
   DFF_X1 \result_reg[7]  (.D(n_171), .CK(n_0), .Q(result[7]), .QN());
   DFF_X1 \result_reg[6]  (.D(n_170), .CK(n_0), .Q(result[6]), .QN());
   DFF_X1 \result_reg[5]  (.D(n_169), .CK(n_0), .Q(result[5]), .QN());
   DFF_X1 \result_reg[4]  (.D(n_168), .CK(n_0), .Q(result[4]), .QN());
   DFF_X1 \result_reg[3]  (.D(n_167), .CK(n_0), .Q(result[3]), .QN());
   DFF_X1 \result_reg[2]  (.D(n_166), .CK(n_0), .Q(result[2]), .QN());
   DFF_X1 \result_reg[1]  (.D(n_165), .CK(n_0), .Q(result[1]), .QN());
   DFF_X1 \result_reg[0]  (.D(n_164), .CK(n_0), .Q(result[0]), .QN());
   CLKGATETST_X1 clk_gate_counter_reg (.CK(clk), .E(en), .SE(1'b0), .GCK(n_1));
   DFF_X1 \counter_reg[5]  (.D(n_233), .CK(n_1), .Q(counter[5]), .QN());
   DFF_X1 \counter_reg[4]  (.D(n_232), .CK(n_1), .Q(counter[4]), .QN());
   DFF_X1 \counter_reg[3]  (.D(n_231), .CK(n_1), .Q(counter[3]), .QN());
   DFF_X1 \counter_reg[2]  (.D(n_230), .CK(n_1), .Q(counter[2]), .QN());
   DFF_X1 \counter_reg[1]  (.D(n_229), .CK(n_1), .Q(counter[1]), .QN());
   DFF_X1 \counter_reg[0]  (.D(n_228), .CK(n_1), .Q(counter[0]), .QN());
   DFF_X1 resetReg_reg (.D(n_162), .CK(clk), .Q(resetReg), .QN());
   MUX2_X1 resetReg_reg_enable_mux_0 (.A(resetReg), .B(n_163), .S(n_335), 
      .Z(n_162));
   CLKGATETST_X1 clk_gate_res_reg (.CK(clk), .E(n_332), .SE(1'b0), .GCK(n_2));
   DFF_X1 \res_reg[64]  (.D(n_298), .CK(n_2), .Q(res[64]), .QN());
   DFF_X1 \res_reg[63]  (.D(n_297), .CK(n_2), .Q(res[63]), .QN());
   DFF_X1 \res_reg[62]  (.D(n_296), .CK(n_2), .Q(res[62]), .QN());
   DFF_X1 \res_reg[61]  (.D(n_295), .CK(n_2), .Q(res[61]), .QN());
   DFF_X1 \res_reg[60]  (.D(n_294), .CK(n_2), .Q(res[60]), .QN());
   DFF_X1 \res_reg[59]  (.D(n_293), .CK(n_2), .Q(res[59]), .QN());
   DFF_X1 \res_reg[58]  (.D(n_292), .CK(n_2), .Q(res[58]), .QN());
   DFF_X1 \res_reg[57]  (.D(n_291), .CK(n_2), .Q(res[57]), .QN());
   DFF_X1 \res_reg[56]  (.D(n_290), .CK(n_2), .Q(res[56]), .QN());
   DFF_X1 \res_reg[55]  (.D(n_289), .CK(n_2), .Q(res[55]), .QN());
   DFF_X1 \res_reg[54]  (.D(n_288), .CK(n_2), .Q(res[54]), .QN());
   DFF_X1 \res_reg[53]  (.D(n_287), .CK(n_2), .Q(res[53]), .QN());
   DFF_X1 \res_reg[52]  (.D(n_286), .CK(n_2), .Q(res[52]), .QN());
   DFF_X1 \res_reg[51]  (.D(n_285), .CK(n_2), .Q(res[51]), .QN());
   DFF_X1 \res_reg[50]  (.D(n_284), .CK(n_2), .Q(res[50]), .QN());
   DFF_X1 \res_reg[49]  (.D(n_283), .CK(n_2), .Q(res[49]), .QN());
   DFF_X1 \res_reg[48]  (.D(n_282), .CK(n_2), .Q(res[48]), .QN());
   DFF_X1 \res_reg[47]  (.D(n_281), .CK(n_2), .Q(res[47]), .QN());
   DFF_X1 \res_reg[46]  (.D(n_280), .CK(n_2), .Q(res[46]), .QN());
   DFF_X1 \res_reg[45]  (.D(n_279), .CK(n_2), .Q(res[45]), .QN());
   DFF_X1 \res_reg[44]  (.D(n_278), .CK(n_2), .Q(res[44]), .QN());
   DFF_X1 \res_reg[43]  (.D(n_277), .CK(n_2), .Q(res[43]), .QN());
   DFF_X1 \res_reg[42]  (.D(n_276), .CK(n_2), .Q(res[42]), .QN());
   DFF_X1 \res_reg[41]  (.D(n_275), .CK(n_2), .Q(res[41]), .QN());
   DFF_X1 \res_reg[40]  (.D(n_274), .CK(n_2), .Q(res[40]), .QN());
   DFF_X1 \res_reg[39]  (.D(n_273), .CK(n_2), .Q(res[39]), .QN());
   DFF_X1 \res_reg[38]  (.D(n_272), .CK(n_2), .Q(res[38]), .QN());
   DFF_X1 \res_reg[37]  (.D(n_271), .CK(n_2), .Q(res[37]), .QN());
   DFF_X1 \res_reg[36]  (.D(n_270), .CK(n_2), .Q(res[36]), .QN());
   DFF_X1 \res_reg[35]  (.D(n_269), .CK(n_2), .Q(res[35]), .QN());
   DFF_X1 \res_reg[34]  (.D(n_268), .CK(n_2), .Q(res[34]), .QN());
   DFF_X1 \res_reg[33]  (.D(n_267), .CK(n_2), .Q(res[33]), .QN());
   DFF_X1 \res_reg[32]  (.D(n_266), .CK(n_2), .Q(res[32]), .QN());
   DFF_X1 \res_reg[31]  (.D(n_265), .CK(n_2), .Q(res[31]), .QN());
   DFF_X1 \res_reg[30]  (.D(n_264), .CK(n_2), .Q(res[30]), .QN());
   DFF_X1 \res_reg[29]  (.D(n_263), .CK(n_2), .Q(res[29]), .QN());
   DFF_X1 \res_reg[28]  (.D(n_262), .CK(n_2), .Q(res[28]), .QN());
   DFF_X1 \res_reg[27]  (.D(n_261), .CK(n_2), .Q(res[27]), .QN());
   DFF_X1 \res_reg[26]  (.D(n_260), .CK(n_2), .Q(res[26]), .QN());
   DFF_X1 \res_reg[25]  (.D(n_259), .CK(n_2), .Q(res[25]), .QN());
   DFF_X1 \res_reg[24]  (.D(n_258), .CK(n_2), .Q(res[24]), .QN());
   DFF_X1 \res_reg[23]  (.D(n_257), .CK(n_2), .Q(res[23]), .QN());
   DFF_X1 \res_reg[22]  (.D(n_256), .CK(n_2), .Q(res[22]), .QN());
   DFF_X1 \res_reg[21]  (.D(n_255), .CK(n_2), .Q(res[21]), .QN());
   DFF_X1 \res_reg[20]  (.D(n_254), .CK(n_2), .Q(res[20]), .QN());
   DFF_X1 \res_reg[19]  (.D(n_253), .CK(n_2), .Q(res[19]), .QN());
   DFF_X1 \res_reg[18]  (.D(n_252), .CK(n_2), .Q(res[18]), .QN());
   DFF_X1 \res_reg[17]  (.D(n_251), .CK(n_2), .Q(res[17]), .QN());
   DFF_X1 \res_reg[16]  (.D(n_250), .CK(n_2), .Q(res[16]), .QN());
   DFF_X1 \res_reg[15]  (.D(n_249), .CK(n_2), .Q(res[15]), .QN());
   DFF_X1 \res_reg[14]  (.D(n_248), .CK(n_2), .Q(res[14]), .QN());
   DFF_X1 \res_reg[13]  (.D(n_247), .CK(n_2), .Q(res[13]), .QN());
   DFF_X1 \res_reg[12]  (.D(n_246), .CK(n_2), .Q(res[12]), .QN());
   DFF_X1 \res_reg[11]  (.D(n_245), .CK(n_2), .Q(res[11]), .QN());
   DFF_X1 \res_reg[10]  (.D(n_244), .CK(n_2), .Q(res[10]), .QN());
   DFF_X1 \res_reg[9]  (.D(n_243), .CK(n_2), .Q(res[9]), .QN());
   DFF_X1 \res_reg[8]  (.D(n_242), .CK(n_2), .Q(res[8]), .QN());
   DFF_X1 \res_reg[7]  (.D(n_241), .CK(n_2), .Q(res[7]), .QN());
   DFF_X1 \res_reg[6]  (.D(n_240), .CK(n_2), .Q(res[6]), .QN());
   DFF_X1 \res_reg[5]  (.D(n_239), .CK(n_2), .Q(res[5]), .QN());
   DFF_X1 \res_reg[4]  (.D(n_238), .CK(n_2), .Q(res[4]), .QN());
   DFF_X1 \res_reg[3]  (.D(n_237), .CK(n_2), .Q(res[3]), .QN());
   DFF_X1 \res_reg[2]  (.D(n_236), .CK(n_2), .Q(res[2]), .QN());
   DFF_X1 \res_reg[1]  (.D(n_235), .CK(n_2), .Q(res[1]), .QN());
   DFF_X1 \res_reg[0]  (.D(n_234), .CK(n_2), .Q(res[0]), .QN());
   HA_X1 i_1_0 (.A(counter[1]), .B(counter[0]), .CO(n_1_0), .S(n_1_3));
   HA_X1 i_1_1 (.A(counter[2]), .B(n_1_0), .CO(n_1_1), .S(n_1_4));
   HA_X1 i_1_2 (.A(counter[3]), .B(n_1_1), .CO(n_1_2), .S(n_1_5));
   HA_X1 i_1_3 (.A(counter[4]), .B(n_1_2), .CO(n_1_7), .S(n_1_6));
   AND2_X1 i_1_4 (.A1(en), .A2(reset), .ZN(n_163));
   AND2_X1 i_1_5 (.A1(n_1_184), .A2(res[1]), .ZN(n_164));
   INV_X1 i_1_6 (.A(n_1_8), .ZN(n_165));
   AOI22_X1 i_1_7 (.A1(res[2]), .A2(n_1_72), .B1(n_1_71), .B2(n_98), .ZN(n_1_8));
   INV_X1 i_1_8 (.A(n_1_9), .ZN(n_166));
   AOI22_X1 i_1_9 (.A1(res[3]), .A2(n_1_72), .B1(n_1_71), .B2(n_99), .ZN(n_1_9));
   INV_X1 i_1_10 (.A(n_1_10), .ZN(n_167));
   AOI22_X1 i_1_11 (.A1(res[4]), .A2(n_1_72), .B1(n_1_71), .B2(n_100), .ZN(
      n_1_10));
   INV_X1 i_1_12 (.A(n_1_11), .ZN(n_168));
   AOI22_X1 i_1_13 (.A1(res[5]), .A2(n_1_72), .B1(n_1_71), .B2(n_101), .ZN(
      n_1_11));
   INV_X1 i_1_14 (.A(n_1_12), .ZN(n_169));
   AOI22_X1 i_1_15 (.A1(res[6]), .A2(n_1_72), .B1(n_1_71), .B2(n_102), .ZN(
      n_1_12));
   INV_X1 i_1_16 (.A(n_1_13), .ZN(n_170));
   AOI22_X1 i_1_17 (.A1(res[7]), .A2(n_1_72), .B1(n_1_71), .B2(n_103), .ZN(
      n_1_13));
   INV_X1 i_1_18 (.A(n_1_14), .ZN(n_171));
   AOI22_X1 i_1_19 (.A1(res[8]), .A2(n_1_72), .B1(n_1_71), .B2(n_104), .ZN(
      n_1_14));
   INV_X1 i_1_20 (.A(n_1_15), .ZN(n_172));
   AOI22_X1 i_1_21 (.A1(res[9]), .A2(n_1_72), .B1(n_1_71), .B2(n_105), .ZN(
      n_1_15));
   INV_X1 i_1_22 (.A(n_1_16), .ZN(n_173));
   AOI22_X1 i_1_23 (.A1(res[10]), .A2(n_1_72), .B1(n_1_71), .B2(n_106), .ZN(
      n_1_16));
   INV_X1 i_1_24 (.A(n_1_17), .ZN(n_174));
   AOI22_X1 i_1_25 (.A1(res[11]), .A2(n_1_72), .B1(n_1_71), .B2(n_107), .ZN(
      n_1_17));
   INV_X1 i_1_26 (.A(n_1_18), .ZN(n_175));
   AOI22_X1 i_1_27 (.A1(res[12]), .A2(n_1_72), .B1(n_1_71), .B2(n_108), .ZN(
      n_1_18));
   INV_X1 i_1_28 (.A(n_1_19), .ZN(n_176));
   AOI22_X1 i_1_29 (.A1(res[13]), .A2(n_1_72), .B1(n_1_71), .B2(n_109), .ZN(
      n_1_19));
   INV_X1 i_1_30 (.A(n_1_20), .ZN(n_177));
   AOI22_X1 i_1_31 (.A1(res[14]), .A2(n_1_72), .B1(n_1_71), .B2(n_110), .ZN(
      n_1_20));
   INV_X1 i_1_32 (.A(n_1_21), .ZN(n_178));
   AOI22_X1 i_1_33 (.A1(res[15]), .A2(n_1_72), .B1(n_1_71), .B2(n_111), .ZN(
      n_1_21));
   INV_X1 i_1_34 (.A(n_1_22), .ZN(n_179));
   AOI22_X1 i_1_35 (.A1(res[16]), .A2(n_1_72), .B1(n_1_71), .B2(n_112), .ZN(
      n_1_22));
   INV_X1 i_1_36 (.A(n_1_23), .ZN(n_180));
   AOI22_X1 i_1_37 (.A1(res[17]), .A2(n_1_72), .B1(n_1_71), .B2(n_113), .ZN(
      n_1_23));
   INV_X1 i_1_38 (.A(n_1_24), .ZN(n_181));
   AOI22_X1 i_1_39 (.A1(res[18]), .A2(n_1_72), .B1(n_1_71), .B2(n_114), .ZN(
      n_1_24));
   INV_X1 i_1_40 (.A(n_1_25), .ZN(n_182));
   AOI22_X1 i_1_41 (.A1(res[19]), .A2(n_1_72), .B1(n_1_71), .B2(n_115), .ZN(
      n_1_25));
   INV_X1 i_1_42 (.A(n_1_26), .ZN(n_183));
   AOI22_X1 i_1_43 (.A1(res[20]), .A2(n_1_72), .B1(n_1_71), .B2(n_116), .ZN(
      n_1_26));
   INV_X1 i_1_44 (.A(n_1_27), .ZN(n_184));
   AOI22_X1 i_1_45 (.A1(res[21]), .A2(n_1_72), .B1(n_1_71), .B2(n_117), .ZN(
      n_1_27));
   INV_X1 i_1_46 (.A(n_1_28), .ZN(n_185));
   AOI22_X1 i_1_47 (.A1(res[22]), .A2(n_1_72), .B1(n_1_71), .B2(n_118), .ZN(
      n_1_28));
   INV_X1 i_1_48 (.A(n_1_29), .ZN(n_186));
   AOI22_X1 i_1_49 (.A1(res[23]), .A2(n_1_72), .B1(n_1_71), .B2(n_119), .ZN(
      n_1_29));
   INV_X1 i_1_50 (.A(n_1_30), .ZN(n_187));
   AOI22_X1 i_1_51 (.A1(res[24]), .A2(n_1_72), .B1(n_1_71), .B2(n_120), .ZN(
      n_1_30));
   INV_X1 i_1_52 (.A(n_1_31), .ZN(n_188));
   AOI22_X1 i_1_53 (.A1(res[25]), .A2(n_1_72), .B1(n_1_71), .B2(n_121), .ZN(
      n_1_31));
   INV_X1 i_1_54 (.A(n_1_32), .ZN(n_189));
   AOI22_X1 i_1_55 (.A1(res[26]), .A2(n_1_72), .B1(n_1_71), .B2(n_122), .ZN(
      n_1_32));
   INV_X1 i_1_56 (.A(n_1_33), .ZN(n_190));
   AOI22_X1 i_1_57 (.A1(res[27]), .A2(n_1_72), .B1(n_1_71), .B2(n_123), .ZN(
      n_1_33));
   INV_X1 i_1_58 (.A(n_1_34), .ZN(n_191));
   AOI22_X1 i_1_59 (.A1(res[28]), .A2(n_1_72), .B1(n_1_71), .B2(n_124), .ZN(
      n_1_34));
   INV_X1 i_1_60 (.A(n_1_35), .ZN(n_192));
   AOI22_X1 i_1_61 (.A1(res[29]), .A2(n_1_72), .B1(n_1_71), .B2(n_125), .ZN(
      n_1_35));
   INV_X1 i_1_62 (.A(n_1_36), .ZN(n_193));
   AOI22_X1 i_1_63 (.A1(res[30]), .A2(n_1_72), .B1(n_1_71), .B2(n_126), .ZN(
      n_1_36));
   INV_X1 i_1_64 (.A(n_1_37), .ZN(n_194));
   AOI22_X1 i_1_65 (.A1(res[31]), .A2(n_1_72), .B1(n_1_71), .B2(n_127), .ZN(
      n_1_37));
   INV_X1 i_1_66 (.A(n_1_38), .ZN(n_195));
   AOI22_X1 i_1_67 (.A1(n_299), .A2(n_1_72), .B1(n_1_71), .B2(n_128), .ZN(n_1_38));
   INV_X1 i_1_68 (.A(n_1_39), .ZN(n_196));
   AOI22_X1 i_1_69 (.A1(n_300), .A2(n_1_72), .B1(n_1_71), .B2(n_129), .ZN(n_1_39));
   INV_X1 i_1_70 (.A(n_1_40), .ZN(n_197));
   AOI22_X1 i_1_71 (.A1(n_301), .A2(n_1_72), .B1(n_1_71), .B2(n_130), .ZN(n_1_40));
   INV_X1 i_1_72 (.A(n_1_41), .ZN(n_198));
   AOI22_X1 i_1_73 (.A1(n_302), .A2(n_1_72), .B1(n_1_71), .B2(n_131), .ZN(n_1_41));
   INV_X1 i_1_74 (.A(n_1_42), .ZN(n_199));
   AOI22_X1 i_1_75 (.A1(n_303), .A2(n_1_72), .B1(n_1_71), .B2(n_132), .ZN(n_1_42));
   INV_X1 i_1_76 (.A(n_1_43), .ZN(n_200));
   AOI22_X1 i_1_77 (.A1(n_304), .A2(n_1_72), .B1(n_1_71), .B2(n_133), .ZN(n_1_43));
   INV_X1 i_1_78 (.A(n_1_44), .ZN(n_201));
   AOI22_X1 i_1_79 (.A1(n_305), .A2(n_1_72), .B1(n_1_71), .B2(n_134), .ZN(n_1_44));
   INV_X1 i_1_80 (.A(n_1_45), .ZN(n_202));
   AOI22_X1 i_1_81 (.A1(n_306), .A2(n_1_72), .B1(n_1_71), .B2(n_135), .ZN(n_1_45));
   INV_X1 i_1_82 (.A(n_1_46), .ZN(n_203));
   AOI22_X1 i_1_83 (.A1(n_307), .A2(n_1_72), .B1(n_1_71), .B2(n_136), .ZN(n_1_46));
   INV_X1 i_1_84 (.A(n_1_47), .ZN(n_204));
   AOI22_X1 i_1_85 (.A1(n_308), .A2(n_1_72), .B1(n_1_71), .B2(n_137), .ZN(n_1_47));
   INV_X1 i_1_86 (.A(n_1_48), .ZN(n_205));
   AOI22_X1 i_1_87 (.A1(n_309), .A2(n_1_72), .B1(n_1_71), .B2(n_138), .ZN(n_1_48));
   INV_X1 i_1_88 (.A(n_1_49), .ZN(n_206));
   AOI22_X1 i_1_89 (.A1(n_310), .A2(n_1_72), .B1(n_1_71), .B2(n_139), .ZN(n_1_49));
   INV_X1 i_1_90 (.A(n_1_50), .ZN(n_207));
   AOI22_X1 i_1_91 (.A1(n_311), .A2(n_1_72), .B1(n_1_71), .B2(n_140), .ZN(n_1_50));
   INV_X1 i_1_92 (.A(n_1_51), .ZN(n_208));
   AOI22_X1 i_1_93 (.A1(n_312), .A2(n_1_72), .B1(n_1_71), .B2(n_141), .ZN(n_1_51));
   INV_X1 i_1_94 (.A(n_1_52), .ZN(n_209));
   AOI22_X1 i_1_95 (.A1(n_313), .A2(n_1_72), .B1(n_1_71), .B2(n_142), .ZN(n_1_52));
   INV_X1 i_1_96 (.A(n_1_53), .ZN(n_210));
   AOI22_X1 i_1_97 (.A1(n_314), .A2(n_1_72), .B1(n_1_71), .B2(n_143), .ZN(n_1_53));
   INV_X1 i_1_98 (.A(n_1_54), .ZN(n_211));
   AOI22_X1 i_1_99 (.A1(n_315), .A2(n_1_72), .B1(n_1_71), .B2(n_144), .ZN(n_1_54));
   INV_X1 i_1_100 (.A(n_1_55), .ZN(n_212));
   AOI22_X1 i_1_101 (.A1(n_316), .A2(n_1_72), .B1(n_1_71), .B2(n_145), .ZN(
      n_1_55));
   INV_X1 i_1_102 (.A(n_1_56), .ZN(n_213));
   AOI22_X1 i_1_103 (.A1(n_317), .A2(n_1_72), .B1(n_1_71), .B2(n_146), .ZN(
      n_1_56));
   INV_X1 i_1_104 (.A(n_1_57), .ZN(n_214));
   AOI22_X1 i_1_105 (.A1(n_318), .A2(n_1_72), .B1(n_1_71), .B2(n_147), .ZN(
      n_1_57));
   INV_X1 i_1_106 (.A(n_1_58), .ZN(n_215));
   AOI22_X1 i_1_107 (.A1(n_319), .A2(n_1_72), .B1(n_1_71), .B2(n_148), .ZN(
      n_1_58));
   INV_X1 i_1_108 (.A(n_1_59), .ZN(n_216));
   AOI22_X1 i_1_109 (.A1(n_320), .A2(n_1_72), .B1(n_1_71), .B2(n_149), .ZN(
      n_1_59));
   INV_X1 i_1_110 (.A(n_1_60), .ZN(n_217));
   AOI22_X1 i_1_111 (.A1(n_321), .A2(n_1_72), .B1(n_1_71), .B2(n_150), .ZN(
      n_1_60));
   INV_X1 i_1_112 (.A(n_1_61), .ZN(n_218));
   AOI22_X1 i_1_113 (.A1(n_322), .A2(n_1_72), .B1(n_1_71), .B2(n_151), .ZN(
      n_1_61));
   INV_X1 i_1_114 (.A(n_1_62), .ZN(n_219));
   AOI22_X1 i_1_115 (.A1(n_323), .A2(n_1_72), .B1(n_1_71), .B2(n_152), .ZN(
      n_1_62));
   INV_X1 i_1_116 (.A(n_1_63), .ZN(n_220));
   AOI22_X1 i_1_117 (.A1(n_324), .A2(n_1_72), .B1(n_1_71), .B2(n_153), .ZN(
      n_1_63));
   INV_X1 i_1_118 (.A(n_1_64), .ZN(n_221));
   AOI22_X1 i_1_119 (.A1(n_325), .A2(n_1_72), .B1(n_1_71), .B2(n_154), .ZN(
      n_1_64));
   INV_X1 i_1_120 (.A(n_1_65), .ZN(n_222));
   AOI22_X1 i_1_121 (.A1(n_326), .A2(n_1_72), .B1(n_1_71), .B2(n_155), .ZN(
      n_1_65));
   INV_X1 i_1_122 (.A(n_1_66), .ZN(n_223));
   AOI22_X1 i_1_123 (.A1(n_327), .A2(n_1_72), .B1(n_1_71), .B2(n_156), .ZN(
      n_1_66));
   INV_X1 i_1_124 (.A(n_1_67), .ZN(n_224));
   AOI22_X1 i_1_125 (.A1(n_328), .A2(n_1_72), .B1(n_1_71), .B2(n_157), .ZN(
      n_1_67));
   INV_X1 i_1_126 (.A(n_1_68), .ZN(n_225));
   AOI22_X1 i_1_127 (.A1(n_329), .A2(n_1_72), .B1(n_1_71), .B2(n_158), .ZN(
      n_1_68));
   INV_X1 i_1_128 (.A(n_1_69), .ZN(n_226));
   AOI22_X1 i_1_129 (.A1(n_330), .A2(n_1_72), .B1(n_1_71), .B2(n_159), .ZN(
      n_1_69));
   INV_X1 i_1_130 (.A(n_1_70), .ZN(n_227));
   AOI22_X1 i_1_131 (.A1(n_331), .A2(n_1_72), .B1(n_1_71), .B2(n_160), .ZN(
      n_1_70));
   NOR2_X1 i_1_132 (.A1(n_335), .A2(n_1_175), .ZN(n_1_71));
   AND2_X1 i_1_133 (.A1(n_1_175), .A2(n_1_184), .ZN(n_1_72));
   AOI211_X1 i_1_134 (.A(counter[0]), .B(n_335), .C1(n_1_186), .C2(counter[5]), 
      .ZN(n_228));
   AND2_X1 i_1_135 (.A1(n_1_73), .A2(n_1_3), .ZN(n_229));
   AND2_X1 i_1_136 (.A1(n_1_73), .A2(n_1_4), .ZN(n_230));
   AND2_X1 i_1_137 (.A1(n_1_73), .A2(n_1_5), .ZN(n_231));
   AND2_X1 i_1_138 (.A1(n_1_73), .A2(n_1_6), .ZN(n_232));
   AND2_X1 i_1_139 (.A1(n_1_178), .A2(n_1_73), .ZN(n_233));
   OAI22_X1 i_1_140 (.A1(en), .A2(counter[5]), .B1(n_335), .B2(n_1_183), 
      .ZN(n_1_73));
   INV_X1 i_1_141 (.A(n_1_74), .ZN(n_234));
   AOI222_X1 i_1_142 (.A1(res[1]), .A2(n_1_180), .B1(n_1_135), .B2(n_3), 
      .C1(in2[1]), .C2(n_1_132), .ZN(n_1_74));
   NAND2_X1 i_1_143 (.A1(n_1_75), .A2(n_1_76), .ZN(n_235));
   AOI22_X1 i_1_144 (.A1(n_4), .A2(n_1_135), .B1(n_1_132), .B2(in2[2]), .ZN(
      n_1_75));
   AOI22_X1 i_1_145 (.A1(res[2]), .A2(n_1_173), .B1(n_1_172), .B2(n_98), 
      .ZN(n_1_76));
   NAND2_X1 i_1_146 (.A1(n_1_77), .A2(n_1_78), .ZN(n_236));
   AOI22_X1 i_1_147 (.A1(n_5), .A2(n_1_135), .B1(n_1_132), .B2(in2[3]), .ZN(
      n_1_77));
   AOI22_X1 i_1_148 (.A1(res[3]), .A2(n_1_173), .B1(n_1_172), .B2(n_99), 
      .ZN(n_1_78));
   NAND2_X1 i_1_149 (.A1(n_1_79), .A2(n_1_80), .ZN(n_237));
   AOI22_X1 i_1_150 (.A1(n_6), .A2(n_1_135), .B1(n_1_132), .B2(in2[4]), .ZN(
      n_1_79));
   AOI22_X1 i_1_151 (.A1(res[4]), .A2(n_1_173), .B1(n_1_172), .B2(n_100), 
      .ZN(n_1_80));
   NAND2_X1 i_1_152 (.A1(n_1_81), .A2(n_1_82), .ZN(n_238));
   AOI22_X1 i_1_153 (.A1(n_7), .A2(n_1_135), .B1(n_1_132), .B2(in2[5]), .ZN(
      n_1_81));
   NAND2_X1 i_1_154 (.A1(n_1_83), .A2(n_1_84), .ZN(n_239));
   AOI22_X1 i_1_155 (.A1(n_8), .A2(n_1_135), .B1(n_1_132), .B2(in2[6]), .ZN(
      n_1_83));
   AOI22_X1 i_1_156 (.A1(res[6]), .A2(n_1_173), .B1(n_1_172), .B2(n_102), 
      .ZN(n_1_84));
   NAND2_X1 i_1_158 (.A1(n_1_85), .A2(n_1_86), .ZN(n_240));
   AOI22_X1 i_1_159 (.A1(n_9), .A2(n_1_135), .B1(n_1_132), .B2(in2[7]), .ZN(
      n_1_85));
   AOI22_X1 i_1_160 (.A1(res[7]), .A2(n_1_173), .B1(n_1_172), .B2(n_103), 
      .ZN(n_1_86));
   NAND2_X1 i_1_161 (.A1(n_1_87), .A2(n_1_88), .ZN(n_241));
   AOI22_X1 i_1_162 (.A1(n_10), .A2(n_1_135), .B1(n_1_132), .B2(in2[8]), 
      .ZN(n_1_87));
   AOI22_X1 i_1_163 (.A1(res[8]), .A2(n_1_173), .B1(n_1_172), .B2(n_104), 
      .ZN(n_1_88));
   NAND2_X1 i_1_164 (.A1(n_1_89), .A2(n_1_90), .ZN(n_242));
   AOI22_X1 i_1_165 (.A1(n_11), .A2(n_1_135), .B1(n_1_132), .B2(in2[9]), 
      .ZN(n_1_89));
   AOI22_X1 i_1_166 (.A1(res[9]), .A2(n_1_173), .B1(n_1_172), .B2(n_105), 
      .ZN(n_1_90));
   NAND2_X1 i_1_167 (.A1(n_1_91), .A2(n_1_92), .ZN(n_243));
   AOI22_X1 i_1_168 (.A1(n_12), .A2(n_1_135), .B1(n_1_132), .B2(in2[10]), 
      .ZN(n_1_91));
   AOI22_X1 i_1_169 (.A1(res[10]), .A2(n_1_173), .B1(n_1_172), .B2(n_106), 
      .ZN(n_1_92));
   NAND2_X1 i_1_170 (.A1(n_1_93), .A2(n_1_94), .ZN(n_244));
   AOI22_X1 i_1_171 (.A1(n_13), .A2(n_1_135), .B1(n_1_132), .B2(in2[11]), 
      .ZN(n_1_93));
   AOI22_X1 i_1_172 (.A1(res[11]), .A2(n_1_173), .B1(n_1_172), .B2(n_107), 
      .ZN(n_1_94));
   NAND2_X1 i_1_173 (.A1(n_1_95), .A2(n_1_96), .ZN(n_245));
   AOI22_X1 i_1_174 (.A1(n_14), .A2(n_1_135), .B1(n_1_132), .B2(in2[12]), 
      .ZN(n_1_95));
   AOI22_X1 i_1_175 (.A1(res[12]), .A2(n_1_173), .B1(n_1_172), .B2(n_108), 
      .ZN(n_1_96));
   NAND2_X1 i_1_176 (.A1(n_1_97), .A2(n_1_98), .ZN(n_246));
   AOI22_X1 i_1_177 (.A1(n_15), .A2(n_1_135), .B1(n_1_132), .B2(in2[13]), 
      .ZN(n_1_97));
   AOI22_X1 i_1_178 (.A1(res[13]), .A2(n_1_173), .B1(n_1_172), .B2(n_109), 
      .ZN(n_1_98));
   NAND2_X1 i_1_179 (.A1(n_1_99), .A2(n_1_100), .ZN(n_247));
   AOI22_X1 i_1_180 (.A1(n_16), .A2(n_1_135), .B1(n_1_132), .B2(in2[14]), 
      .ZN(n_1_99));
   AOI22_X1 i_1_181 (.A1(res[14]), .A2(n_1_173), .B1(n_1_172), .B2(n_110), 
      .ZN(n_1_100));
   NAND2_X1 i_1_182 (.A1(n_1_101), .A2(n_1_102), .ZN(n_248));
   AOI22_X1 i_1_183 (.A1(n_17), .A2(n_1_135), .B1(n_1_132), .B2(in2[15]), 
      .ZN(n_1_101));
   AOI22_X1 i_1_184 (.A1(res[15]), .A2(n_1_173), .B1(n_1_172), .B2(n_111), 
      .ZN(n_1_102));
   NAND2_X1 i_1_185 (.A1(n_1_103), .A2(n_1_104), .ZN(n_249));
   AOI22_X1 i_1_186 (.A1(n_18), .A2(n_1_135), .B1(n_1_132), .B2(in2[16]), 
      .ZN(n_1_103));
   AOI22_X1 i_1_187 (.A1(res[16]), .A2(n_1_173), .B1(n_1_172), .B2(n_112), 
      .ZN(n_1_104));
   NAND2_X1 i_1_188 (.A1(n_1_105), .A2(n_1_106), .ZN(n_250));
   AOI22_X1 i_1_189 (.A1(n_19), .A2(n_1_135), .B1(n_1_132), .B2(in2[17]), 
      .ZN(n_1_105));
   AOI22_X1 i_1_190 (.A1(res[17]), .A2(n_1_173), .B1(n_1_172), .B2(n_113), 
      .ZN(n_1_106));
   NAND2_X1 i_1_191 (.A1(n_1_107), .A2(n_1_108), .ZN(n_251));
   AOI22_X1 i_1_192 (.A1(n_20), .A2(n_1_135), .B1(n_1_132), .B2(in2[18]), 
      .ZN(n_1_107));
   AOI22_X1 i_1_193 (.A1(res[18]), .A2(n_1_173), .B1(n_1_172), .B2(n_114), 
      .ZN(n_1_108));
   NAND2_X1 i_1_194 (.A1(n_1_109), .A2(n_1_110), .ZN(n_252));
   AOI22_X1 i_1_195 (.A1(n_21), .A2(n_1_135), .B1(n_1_132), .B2(in2[19]), 
      .ZN(n_1_109));
   AOI22_X1 i_1_196 (.A1(res[19]), .A2(n_1_173), .B1(n_1_172), .B2(n_115), 
      .ZN(n_1_110));
   NAND2_X1 i_1_197 (.A1(n_1_111), .A2(n_1_112), .ZN(n_253));
   AOI22_X1 i_1_198 (.A1(n_22), .A2(n_1_135), .B1(n_1_132), .B2(in2[20]), 
      .ZN(n_1_111));
   AOI22_X1 i_1_199 (.A1(res[20]), .A2(n_1_173), .B1(n_1_172), .B2(n_116), 
      .ZN(n_1_112));
   NAND2_X1 i_1_200 (.A1(n_1_113), .A2(n_1_114), .ZN(n_254));
   AOI22_X1 i_1_201 (.A1(n_23), .A2(n_1_135), .B1(n_1_132), .B2(in2[21]), 
      .ZN(n_1_113));
   AOI22_X1 i_1_202 (.A1(res[21]), .A2(n_1_173), .B1(n_1_172), .B2(n_117), 
      .ZN(n_1_114));
   NAND2_X1 i_1_203 (.A1(n_1_115), .A2(n_1_116), .ZN(n_255));
   AOI22_X1 i_1_204 (.A1(n_24), .A2(n_1_135), .B1(n_1_132), .B2(in2[22]), 
      .ZN(n_1_115));
   AOI22_X1 i_1_205 (.A1(res[22]), .A2(n_1_173), .B1(n_1_172), .B2(n_118), 
      .ZN(n_1_116));
   NAND2_X1 i_1_206 (.A1(n_1_117), .A2(n_1_118), .ZN(n_256));
   AOI22_X1 i_1_207 (.A1(n_25), .A2(n_1_135), .B1(n_1_132), .B2(in2[23]), 
      .ZN(n_1_117));
   AOI22_X1 i_1_208 (.A1(res[23]), .A2(n_1_173), .B1(n_1_172), .B2(n_119), 
      .ZN(n_1_118));
   NAND2_X1 i_1_209 (.A1(n_1_119), .A2(n_1_120), .ZN(n_257));
   AOI22_X1 i_1_210 (.A1(n_26), .A2(n_1_135), .B1(n_1_132), .B2(in2[24]), 
      .ZN(n_1_119));
   AOI22_X1 i_1_211 (.A1(res[24]), .A2(n_1_173), .B1(n_1_172), .B2(n_120), 
      .ZN(n_1_120));
   NAND2_X1 i_1_212 (.A1(n_1_121), .A2(n_1_122), .ZN(n_258));
   AOI22_X1 i_1_213 (.A1(n_27), .A2(n_1_135), .B1(n_1_132), .B2(in2[25]), 
      .ZN(n_1_121));
   AOI22_X1 i_1_214 (.A1(res[25]), .A2(n_1_173), .B1(n_1_172), .B2(n_121), 
      .ZN(n_1_122));
   NAND2_X1 i_1_215 (.A1(n_1_123), .A2(n_1_124), .ZN(n_259));
   AOI22_X1 i_1_216 (.A1(n_28), .A2(n_1_135), .B1(n_1_132), .B2(in2[26]), 
      .ZN(n_1_123));
   AOI22_X1 i_1_217 (.A1(res[26]), .A2(n_1_173), .B1(n_1_172), .B2(n_122), 
      .ZN(n_1_124));
   NAND2_X1 i_1_218 (.A1(n_1_125), .A2(n_1_126), .ZN(n_260));
   AOI22_X1 i_1_219 (.A1(n_29), .A2(n_1_135), .B1(n_1_132), .B2(in2[27]), 
      .ZN(n_1_125));
   AOI22_X1 i_1_220 (.A1(res[27]), .A2(n_1_173), .B1(n_1_172), .B2(n_123), 
      .ZN(n_1_126));
   NAND2_X1 i_1_221 (.A1(n_1_127), .A2(n_1_128), .ZN(n_261));
   AOI22_X1 i_1_222 (.A1(n_30), .A2(n_1_135), .B1(n_1_132), .B2(in2[28]), 
      .ZN(n_1_127));
   AOI22_X1 i_1_223 (.A1(res[28]), .A2(n_1_173), .B1(n_1_172), .B2(n_124), 
      .ZN(n_1_128));
   NAND2_X1 i_1_224 (.A1(n_1_129), .A2(n_1_130), .ZN(n_262));
   AOI22_X1 i_1_225 (.A1(n_31), .A2(n_1_135), .B1(n_1_132), .B2(in2[29]), 
      .ZN(n_1_129));
   AOI22_X1 i_1_226 (.A1(res[29]), .A2(n_1_173), .B1(n_1_172), .B2(n_125), 
      .ZN(n_1_130));
   NAND2_X1 i_1_227 (.A1(n_1_131), .A2(n_1_133), .ZN(n_263));
   AOI22_X1 i_1_228 (.A1(n_32), .A2(n_1_135), .B1(n_1_132), .B2(in2[30]), 
      .ZN(n_1_131));
   NOR4_X1 i_1_157 (.A1(n_1_182), .A2(in2[31]), .A3(resetReg), .A4(reset), 
      .ZN(n_1_132));
   AOI22_X1 i_1_230 (.A1(res[30]), .A2(n_1_173), .B1(n_1_172), .B2(n_126), 
      .ZN(n_1_133));
   INV_X1 i_1_231 (.A(n_1_134), .ZN(n_264));
   AOI22_X1 i_1_232 (.A1(n_1_180), .A2(n_1_136), .B1(n_1_135), .B2(n_33), 
      .ZN(n_1_134));
   AND2_X1 i_1_229 (.A1(in2[31]), .A2(n_1_170), .ZN(n_1_135));
   MUX2_X1 i_1_234 (.A(res[31]), .B(n_127), .S(n_1_174), .Z(n_1_136));
   INV_X1 i_1_235 (.A(n_1_137), .ZN(n_265));
   AOI222_X1 i_1_236 (.A1(n_128), .A2(n_1_172), .B1(n_1_169), .B2(in1[0]), 
      .C1(n_1_173), .C2(n_299), .ZN(n_1_137));
   INV_X1 i_1_237 (.A(n_1_138), .ZN(n_266));
   AOI222_X1 i_1_238 (.A1(n_1_169), .A2(m[1]), .B1(n_129), .B2(n_1_172), 
      .C1(n_300), .C2(n_1_173), .ZN(n_1_138));
   INV_X1 i_1_239 (.A(n_1_139), .ZN(n_267));
   AOI222_X1 i_1_240 (.A1(n_1_169), .A2(m[2]), .B1(n_130), .B2(n_1_172), 
      .C1(n_301), .C2(n_1_173), .ZN(n_1_139));
   INV_X1 i_1_241 (.A(n_1_140), .ZN(n_268));
   AOI222_X1 i_1_242 (.A1(n_1_169), .A2(m[3]), .B1(n_131), .B2(n_1_172), 
      .C1(n_302), .C2(n_1_173), .ZN(n_1_140));
   INV_X1 i_1_243 (.A(n_1_141), .ZN(n_269));
   AOI222_X1 i_1_244 (.A1(n_1_169), .A2(m[4]), .B1(n_132), .B2(n_1_172), 
      .C1(n_303), .C2(n_1_173), .ZN(n_1_141));
   INV_X1 i_1_245 (.A(n_1_142), .ZN(n_270));
   AOI222_X1 i_1_246 (.A1(n_1_169), .A2(m[5]), .B1(n_133), .B2(n_1_172), 
      .C1(n_304), .C2(n_1_173), .ZN(n_1_142));
   INV_X1 i_1_247 (.A(n_1_143), .ZN(n_271));
   AOI222_X1 i_1_248 (.A1(n_1_169), .A2(m[6]), .B1(n_134), .B2(n_1_172), 
      .C1(n_305), .C2(n_1_173), .ZN(n_1_143));
   INV_X1 i_1_249 (.A(n_1_144), .ZN(n_272));
   AOI222_X1 i_1_250 (.A1(n_1_169), .A2(m[7]), .B1(n_135), .B2(n_1_172), 
      .C1(n_306), .C2(n_1_173), .ZN(n_1_144));
   INV_X1 i_1_251 (.A(n_1_145), .ZN(n_273));
   AOI222_X1 i_1_252 (.A1(n_1_169), .A2(m[8]), .B1(n_136), .B2(n_1_172), 
      .C1(n_307), .C2(n_1_173), .ZN(n_1_145));
   INV_X1 i_1_253 (.A(n_1_146), .ZN(n_274));
   AOI222_X1 i_1_254 (.A1(n_1_169), .A2(m[9]), .B1(n_137), .B2(n_1_172), 
      .C1(n_308), .C2(n_1_173), .ZN(n_1_146));
   INV_X1 i_1_255 (.A(n_1_147), .ZN(n_275));
   AOI222_X1 i_1_256 (.A1(n_1_169), .A2(m[10]), .B1(n_138), .B2(n_1_172), 
      .C1(n_309), .C2(n_1_173), .ZN(n_1_147));
   INV_X1 i_1_257 (.A(n_1_148), .ZN(n_276));
   AOI222_X1 i_1_258 (.A1(n_1_169), .A2(m[11]), .B1(n_139), .B2(n_1_172), 
      .C1(n_310), .C2(n_1_173), .ZN(n_1_148));
   INV_X1 i_1_259 (.A(n_1_149), .ZN(n_277));
   AOI222_X1 i_1_260 (.A1(n_1_169), .A2(m[12]), .B1(n_140), .B2(n_1_172), 
      .C1(n_311), .C2(n_1_173), .ZN(n_1_149));
   INV_X1 i_1_261 (.A(n_1_150), .ZN(n_278));
   AOI222_X1 i_1_262 (.A1(n_1_169), .A2(m[13]), .B1(n_141), .B2(n_1_172), 
      .C1(n_312), .C2(n_1_173), .ZN(n_1_150));
   INV_X1 i_1_263 (.A(n_1_151), .ZN(n_279));
   AOI222_X1 i_1_264 (.A1(n_1_169), .A2(m[14]), .B1(n_142), .B2(n_1_172), 
      .C1(n_313), .C2(n_1_173), .ZN(n_1_151));
   INV_X1 i_1_265 (.A(n_1_152), .ZN(n_280));
   AOI222_X1 i_1_266 (.A1(n_1_169), .A2(m[15]), .B1(n_143), .B2(n_1_172), 
      .C1(n_314), .C2(n_1_173), .ZN(n_1_152));
   INV_X1 i_1_267 (.A(n_1_153), .ZN(n_281));
   AOI222_X1 i_1_268 (.A1(n_1_169), .A2(m[16]), .B1(n_144), .B2(n_1_172), 
      .C1(n_315), .C2(n_1_173), .ZN(n_1_153));
   INV_X1 i_1_269 (.A(n_1_154), .ZN(n_282));
   AOI222_X1 i_1_270 (.A1(n_1_169), .A2(m[17]), .B1(n_145), .B2(n_1_172), 
      .C1(n_316), .C2(n_1_173), .ZN(n_1_154));
   INV_X1 i_1_271 (.A(n_1_155), .ZN(n_283));
   AOI222_X1 i_1_233 (.A1(n_1_169), .A2(m[18]), .B1(n_146), .B2(n_1_172), 
      .C1(n_317), .C2(n_1_173), .ZN(n_1_155));
   INV_X1 i_1_272 (.A(n_1_156), .ZN(n_284));
   AOI222_X1 i_1_273 (.A1(n_1_169), .A2(m[19]), .B1(n_147), .B2(n_1_172), 
      .C1(n_318), .C2(n_1_173), .ZN(n_1_156));
   INV_X1 i_1_275 (.A(n_1_157), .ZN(n_285));
   AOI222_X1 i_1_276 (.A1(n_1_169), .A2(m[20]), .B1(n_148), .B2(n_1_172), 
      .C1(n_319), .C2(n_1_173), .ZN(n_1_157));
   INV_X1 i_1_277 (.A(n_1_158), .ZN(n_286));
   AOI222_X1 i_1_278 (.A1(n_1_169), .A2(m[21]), .B1(n_149), .B2(n_1_172), 
      .C1(n_320), .C2(n_1_173), .ZN(n_1_158));
   INV_X1 i_1_279 (.A(n_1_159), .ZN(n_287));
   AOI222_X1 i_1_280 (.A1(n_1_169), .A2(m[22]), .B1(n_150), .B2(n_1_172), 
      .C1(n_321), .C2(n_1_173), .ZN(n_1_159));
   INV_X1 i_1_281 (.A(n_1_160), .ZN(n_288));
   AOI222_X1 i_1_282 (.A1(n_1_169), .A2(m[23]), .B1(n_151), .B2(n_1_172), 
      .C1(n_322), .C2(n_1_173), .ZN(n_1_160));
   INV_X1 i_1_283 (.A(n_1_161), .ZN(n_289));
   AOI222_X1 i_1_284 (.A1(n_1_169), .A2(m[24]), .B1(n_152), .B2(n_1_172), 
      .C1(n_323), .C2(n_1_173), .ZN(n_1_161));
   INV_X1 i_1_285 (.A(n_1_162), .ZN(n_290));
   AOI222_X1 i_1_286 (.A1(n_1_169), .A2(m[25]), .B1(n_153), .B2(n_1_172), 
      .C1(n_324), .C2(n_1_173), .ZN(n_1_162));
   INV_X1 i_1_287 (.A(n_1_163), .ZN(n_291));
   AOI222_X1 i_1_288 (.A1(n_1_169), .A2(m[26]), .B1(n_154), .B2(n_1_172), 
      .C1(n_325), .C2(n_1_173), .ZN(n_1_163));
   INV_X1 i_1_289 (.A(n_1_164), .ZN(n_292));
   AOI222_X1 i_1_290 (.A1(n_1_169), .A2(m[27]), .B1(n_155), .B2(n_1_172), 
      .C1(n_326), .C2(n_1_173), .ZN(n_1_164));
   INV_X1 i_1_291 (.A(n_1_165), .ZN(n_293));
   AOI222_X1 i_1_292 (.A1(n_1_169), .A2(m[28]), .B1(n_156), .B2(n_1_172), 
      .C1(n_327), .C2(n_1_173), .ZN(n_1_165));
   INV_X1 i_1_293 (.A(n_1_166), .ZN(n_294));
   AOI222_X1 i_1_294 (.A1(n_1_169), .A2(m[29]), .B1(n_157), .B2(n_1_172), 
      .C1(n_328), .C2(n_1_173), .ZN(n_1_166));
   INV_X1 i_1_295 (.A(n_1_167), .ZN(n_295));
   AOI222_X1 i_1_296 (.A1(n_1_169), .A2(m[30]), .B1(n_158), .B2(n_1_172), 
      .C1(n_329), .C2(n_1_173), .ZN(n_1_167));
   INV_X1 i_1_297 (.A(n_1_168), .ZN(n_296));
   AOI222_X1 i_1_298 (.A1(n_159), .A2(n_1_172), .B1(n_1_169), .B2(m[31]), 
      .C1(n_330), .C2(n_1_173), .ZN(n_1_168));
   AND2_X1 i_1_274 (.A1(in2[0]), .A2(n_1_170), .ZN(n_1_169));
   NOR3_X1 i_1_299 (.A1(n_1_182), .A2(resetReg), .A3(reset), .ZN(n_1_170));
   INV_X1 i_1_301 (.A(n_1_171), .ZN(n_297));
   AOI22_X1 i_1_302 (.A1(n_160), .A2(n_1_172), .B1(n_1_173), .B2(n_331), 
      .ZN(n_1_171));
   AND3_X1 i_1_305 (.A1(n_161), .A2(n_1_180), .A3(n_1_174), .ZN(n_298));
   MUX2_X1 i_1_312 (.A(res[32]), .B(n_65), .S(res[0]), .Z(n_299));
   MUX2_X1 i_1_313 (.A(res[33]), .B(n_66), .S(res[0]), .Z(n_300));
   MUX2_X1 i_1_314 (.A(res[34]), .B(n_67), .S(res[0]), .Z(n_301));
   MUX2_X1 i_1_315 (.A(res[35]), .B(n_68), .S(res[0]), .Z(n_302));
   MUX2_X1 i_1_316 (.A(res[36]), .B(n_69), .S(res[0]), .Z(n_303));
   MUX2_X1 i_1_317 (.A(res[37]), .B(n_70), .S(res[0]), .Z(n_304));
   MUX2_X1 i_1_318 (.A(res[38]), .B(n_71), .S(res[0]), .Z(n_305));
   MUX2_X1 i_1_319 (.A(res[39]), .B(n_72), .S(res[0]), .Z(n_306));
   MUX2_X1 i_1_320 (.A(res[40]), .B(n_73), .S(res[0]), .Z(n_307));
   MUX2_X1 i_1_321 (.A(res[41]), .B(n_74), .S(res[0]), .Z(n_308));
   MUX2_X1 i_1_322 (.A(res[42]), .B(n_75), .S(res[0]), .Z(n_309));
   MUX2_X1 i_1_323 (.A(res[43]), .B(n_76), .S(res[0]), .Z(n_310));
   MUX2_X1 i_1_324 (.A(res[44]), .B(n_77), .S(res[0]), .Z(n_311));
   MUX2_X1 i_1_325 (.A(res[45]), .B(n_78), .S(res[0]), .Z(n_312));
   MUX2_X1 i_1_326 (.A(res[46]), .B(n_79), .S(res[0]), .Z(n_313));
   MUX2_X1 i_1_327 (.A(res[47]), .B(n_80), .S(res[0]), .Z(n_314));
   MUX2_X1 i_1_300 (.A(res[48]), .B(n_81), .S(res[0]), .Z(n_315));
   MUX2_X1 i_1_303 (.A(res[49]), .B(n_82), .S(res[0]), .Z(n_316));
   MUX2_X1 i_1_304 (.A(res[50]), .B(n_83), .S(res[0]), .Z(n_317));
   MUX2_X1 i_1_306 (.A(res[51]), .B(n_84), .S(res[0]), .Z(n_318));
   MUX2_X1 i_1_332 (.A(res[52]), .B(n_85), .S(res[0]), .Z(n_319));
   MUX2_X1 i_1_333 (.A(res[53]), .B(n_86), .S(res[0]), .Z(n_320));
   MUX2_X1 i_1_334 (.A(res[54]), .B(n_87), .S(res[0]), .Z(n_321));
   MUX2_X1 i_1_335 (.A(res[55]), .B(n_88), .S(res[0]), .Z(n_322));
   MUX2_X1 i_1_336 (.A(res[56]), .B(n_89), .S(res[0]), .Z(n_323));
   MUX2_X1 i_1_337 (.A(res[57]), .B(n_90), .S(res[0]), .Z(n_324));
   MUX2_X1 i_1_338 (.A(res[58]), .B(n_91), .S(res[0]), .Z(n_325));
   MUX2_X1 i_1_339 (.A(res[59]), .B(n_92), .S(res[0]), .Z(n_326));
   MUX2_X1 i_1_340 (.A(res[60]), .B(n_93), .S(res[0]), .Z(n_327));
   MUX2_X1 i_1_341 (.A(res[61]), .B(n_94), .S(res[0]), .Z(n_328));
   MUX2_X1 i_1_342 (.A(res[62]), .B(n_95), .S(res[0]), .Z(n_329));
   MUX2_X1 i_1_343 (.A(res[63]), .B(n_96), .S(res[0]), .Z(n_330));
   MUX2_X1 i_1_344 (.A(res[64]), .B(n_97), .S(res[0]), .Z(n_331));
   NOR3_X1 i_1_307 (.A1(n_1_188), .A2(reset), .A3(resetReg), .ZN(n_332));
   NAND2_X1 i_1_308 (.A1(n_1_184), .A2(n_1_176), .ZN(n_333));
   AOI21_X1 i_1_309 (.A(n_335), .B1(n_1_176), .B2(en), .ZN(n_334));
   INV_X1 i_1_310 (.A(n_1_184), .ZN(n_335));
   OAI21_X1 i_1_311 (.A(en), .B1(reset), .B2(resetReg), .ZN(n_1_184));
   MUX2_X1 i_1_355 (.A(in1[1]), .B(n_34), .S(in1[31]), .Z(m[1]));
   MUX2_X1 i_1_356 (.A(in1[2]), .B(n_35), .S(in1[31]), .Z(m[2]));
   MUX2_X1 i_1_357 (.A(in1[3]), .B(n_36), .S(in1[31]), .Z(m[3]));
   MUX2_X1 i_1_358 (.A(in1[4]), .B(n_37), .S(in1[31]), .Z(m[4]));
   MUX2_X1 i_1_359 (.A(in1[5]), .B(n_38), .S(in1[31]), .Z(m[5]));
   MUX2_X1 i_1_360 (.A(in1[6]), .B(n_39), .S(in1[31]), .Z(m[6]));
   MUX2_X1 i_1_361 (.A(in1[7]), .B(n_40), .S(in1[31]), .Z(m[7]));
   MUX2_X1 i_1_362 (.A(in1[8]), .B(n_41), .S(in1[31]), .Z(m[8]));
   MUX2_X1 i_1_363 (.A(in1[9]), .B(n_42), .S(in1[31]), .Z(m[9]));
   MUX2_X1 i_1_364 (.A(in1[10]), .B(n_43), .S(in1[31]), .Z(m[10]));
   MUX2_X1 i_1_365 (.A(in1[11]), .B(n_44), .S(in1[31]), .Z(m[11]));
   MUX2_X1 i_1_366 (.A(in1[12]), .B(n_45), .S(in1[31]), .Z(m[12]));
   MUX2_X1 i_1_367 (.A(in1[13]), .B(n_46), .S(in1[31]), .Z(m[13]));
   MUX2_X1 i_1_368 (.A(in1[14]), .B(n_47), .S(in1[31]), .Z(m[14]));
   MUX2_X1 i_1_369 (.A(in1[15]), .B(n_48), .S(in1[31]), .Z(m[15]));
   MUX2_X1 i_1_370 (.A(in1[16]), .B(n_49), .S(in1[31]), .Z(m[16]));
   MUX2_X1 i_1_371 (.A(in1[17]), .B(n_50), .S(in1[31]), .Z(m[17]));
   MUX2_X1 i_1_328 (.A(in1[18]), .B(n_51), .S(in1[31]), .Z(m[18]));
   MUX2_X1 i_1_329 (.A(in1[19]), .B(n_52), .S(in1[31]), .Z(m[19]));
   MUX2_X1 i_1_374 (.A(in1[20]), .B(n_53), .S(in1[31]), .Z(m[20]));
   MUX2_X1 i_1_375 (.A(in1[21]), .B(n_54), .S(in1[31]), .Z(m[21]));
   MUX2_X1 i_1_376 (.A(in1[22]), .B(n_55), .S(in1[31]), .Z(m[22]));
   MUX2_X1 i_1_377 (.A(in1[23]), .B(n_56), .S(in1[31]), .Z(m[23]));
   MUX2_X1 i_1_378 (.A(in1[24]), .B(n_57), .S(in1[31]), .Z(m[24]));
   MUX2_X1 i_1_379 (.A(in1[25]), .B(n_58), .S(in1[31]), .Z(m[25]));
   MUX2_X1 i_1_380 (.A(in1[26]), .B(n_59), .S(in1[31]), .Z(m[26]));
   MUX2_X1 i_1_381 (.A(in1[27]), .B(n_60), .S(in1[31]), .Z(m[27]));
   MUX2_X1 i_1_382 (.A(in1[28]), .B(n_61), .S(in1[31]), .Z(m[28]));
   MUX2_X1 i_1_383 (.A(in1[29]), .B(n_62), .S(in1[31]), .Z(m[29]));
   MUX2_X1 i_1_384 (.A(in1[30]), .B(n_63), .S(in1[31]), .Z(m[30]));
   AND2_X1 i_1_385 (.A1(in1[31]), .A2(n_64), .ZN(m[31]));
   INV_X1 i_1_330 (.A(en), .ZN(n_1_188));
   AOI22_X1 i_1_331 (.A1(res[5]), .A2(n_1_173), .B1(n_101), .B2(n_1_172), 
      .ZN(n_1_82));
   AND2_X1 i_1_345 (.A1(n_1_180), .A2(n_1_174), .ZN(n_1_172));
   NOR2_X1 i_1_346 (.A1(n_1_179), .A2(n_1_174), .ZN(n_1_173));
   NOR2_X1 i_1_347 (.A1(n_1_176), .A2(n_1_175), .ZN(n_1_174));
   XNOR2_X1 i_1_348 (.A(in2[31]), .B(in1[31]), .ZN(n_1_175));
   NAND4_X1 i_1_349 (.A1(counter[0]), .A2(n_1_187), .A3(n_1_177), .A4(n_1_178), 
      .ZN(n_1_176));
   NOR3_X1 i_1_350 (.A1(n_1_5), .A2(n_1_4), .A3(n_1_3), .ZN(n_1_177));
   XOR2_X1 i_1_351 (.A(counter[5]), .B(n_1_7), .Z(n_1_178));
   INV_X1 i_1_352 (.A(n_1_180), .ZN(n_1_179));
   NOR3_X1 i_1_353 (.A1(reset), .A2(resetReg), .A3(n_1_181), .ZN(n_1_180));
   INV_X1 i_1_354 (.A(n_1_182), .ZN(n_1_181));
   OAI21_X1 i_1_372 (.A(n_1_183), .B1(n_1_189), .B2(counter[4]), .ZN(n_1_182));
   NOR2_X1 i_1_373 (.A1(counter[0]), .A2(n_1_185), .ZN(n_1_183));
   INV_X1 i_1_386 (.A(n_1_186), .ZN(n_1_185));
   NOR4_X1 i_1_387 (.A1(counter[4]), .A2(counter[3]), .A3(counter[2]), .A4(
      counter[1]), .ZN(n_1_186));
   INV_X1 i_1_388 (.A(n_1_6), .ZN(n_1_187));
   INV_X1 i_1_389 (.A(counter[5]), .ZN(n_1_189));
endmodule

module registerNbits__0_28(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module integrationMult(inputA, inputB, clk, reset, en, result);
   input [31:0]inputA;
   input [31:0]inputB;
   input clk;
   input reset;
   input en;
   output [63:0]result;

   wire [31:0]A_reg;
   wire [31:0]B_reg;
   wire enableOutput;
   wire [31:0]outB_reg;
   wire [31:0]outA_reg;

   registerNbits__0_22 regA (.clk(clk), .reset(reset), .en(en), .inp(inputA), 
      .out(A_reg));
   registerNbits__0_25 regB (.clk(clk), .reset(reset), .en(en), .inp(inputB), 
      .out(B_reg));
   sequentialmultiplier SM (.in1(A_reg), .in2(B_reg), .clk(clk), .reset(reset), 
      .en(en), .result({outA_reg[31], outA_reg[30], outA_reg[29], outA_reg[28], 
      outA_reg[27], outA_reg[26], outA_reg[25], outA_reg[24], outA_reg[23], 
      outA_reg[22], outA_reg[21], outA_reg[20], outA_reg[19], outA_reg[18], 
      outA_reg[17], outA_reg[16], outA_reg[15], outA_reg[14], outA_reg[13], 
      outA_reg[12], outA_reg[11], outA_reg[10], outA_reg[9], outA_reg[8], 
      outA_reg[7], outA_reg[6], outA_reg[5], outA_reg[4], outA_reg[3], 
      outA_reg[2], outA_reg[1], outA_reg[0], outB_reg[31], outB_reg[30], 
      outB_reg[29], outB_reg[28], outB_reg[27], outB_reg[26], outB_reg[25], 
      outB_reg[24], outB_reg[23], outB_reg[22], outB_reg[21], outB_reg[20], 
      outB_reg[19], outB_reg[18], outB_reg[17], outB_reg[16], outB_reg[15], 
      outB_reg[14], outB_reg[13], outB_reg[12], outB_reg[11], outB_reg[10], 
      outB_reg[9], outB_reg[8], outB_reg[7], outB_reg[6], outB_reg[5], 
      outB_reg[4], outB_reg[3], outB_reg[2], outB_reg[1], outB_reg[0]}), 
      .enableOutput(enableOutput));
   registerNbits__0_28 outB (.clk(clk), .reset(reset), .en(enableOutput), 
      .inp(outA_reg), .out({result[63], result[62], result[61], result[60], 
      result[59], result[58], result[57], result[56], result[55], result[54], 
      result[53], result[52], result[51], result[50], result[49], result[48], 
      result[47], result[46], result[45], result[44], result[43], result[42], 
      result[41], result[40], result[39], result[38], result[37], result[36], 
      result[35], result[34], result[33], result[32]}));
   registerNbits outA (.clk(clk), .reset(reset), .en(enableOutput), .inp(
      outB_reg), .out({result[31], result[30], result[29], result[28], 
      result[27], result[26], result[25], result[24], result[23], result[22], 
      result[21], result[20], result[19], result[18], result[17], result[16], 
      result[15], result[14], result[13], result[12], result[11], result[10], 
      result[9], result[8], result[7], result[6], result[5], result[4], 
      result[3], result[2], result[1], result[0]}));
endmodule
