module RCA8(A,B,cin,cout,sum);
input [7:0]A,B;
input cin;
output [7:0]sum;
output cout;
wire [6:0] carry;

FullAdder FA1 (A[0],B[0],cin,sum[0],carry[0]);
FullAdder FA2 (A[1],B[1],carry[0],sum[1],carry[1]);
FullAdder FA3 (A[2],B[2],carry[1],sum[2],carry[2]);
FullAdder FA4 (A[3],B[3],carry[2],sum[3],carry[3]);
FullAdder FA5 (A[4],B[4],carry[3],sum[4],carry[4]);
FullAdder FA6 (A[5],B[5],carry[4],sum[5],carry[5]);
FullAdder FA7 (A[6],B[6],carry[5],sum[6],carry[6]);
FullAdder FA8 (A[7],B[7],carry[6],sum[7],cout);

endmodule