
// 	Fri Dec 23 14:43:54 2022
//	vlsi
//	localhost.localdomain

module registerNbits (clk_CTS_0_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_2;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid1_3;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_2), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_2), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_2), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_2), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_2), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_2), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_2), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_2), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_2), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_2), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_2), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_2), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_2), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_2), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_2), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_2), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_2), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_2), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_2), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_2), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_2), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_2), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_2), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_2), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_2), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_2), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_2), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_2), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_2), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_2), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_2), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid1_2), .D (n_33));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n_tid1_3), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X3 CTS_L3_c_tid1_3 (.Z (CTS_n_tid1_2), .A (CTS_n_tid1_3));

endmodule //registerNbits

module registerNbits__0_28 (clk_CTS_0_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_2;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid1_3;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_2), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_2), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_2), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_2), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_2), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_2), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_2), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_2), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_2), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_2), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_2), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_2), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_2), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_2), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_2), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_2), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_2), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_2), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_2), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_2), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_2), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_2), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_2), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_2), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_2), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_2), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_2), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_2), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_2), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_2), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_2), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid1_2), .D (n_33));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n_tid1_3), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X3 CTS_L3_c_tid1_3 (.Z (CTS_n_tid1_2), .A (CTS_n_tid1_3));

endmodule //registerNbits__0_28

module datapath__0_11 (p_0, p_1);

output [64:0] p_0;
input [64:0] p_1;
wire n_61;
wire n_0;
wire n_60;
wire n_59;
wire n_58;
wire n_1;
wire n_57;
wire n_56;
wire n_2;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_3;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_4;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_5;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;


INV_X1 i_137 (.ZN (n_73), .A (p_1[63]));
INV_X1 i_136 (.ZN (n_72), .A (p_1[60]));
INV_X1 i_135 (.ZN (n_71), .A (p_1[55]));
INV_X1 i_134 (.ZN (n_70), .A (p_1[51]));
INV_X1 i_133 (.ZN (n_69), .A (p_1[42]));
INV_X1 i_132 (.ZN (n_68), .A (p_1[40]));
INV_X1 i_131 (.ZN (n_67), .A (p_1[36]));
INV_X1 i_130 (.ZN (n_66), .A (p_1[31]));
INV_X1 i_129 (.ZN (n_65), .A (p_1[26]));
INV_X1 i_128 (.ZN (n_64), .A (p_1[21]));
INV_X1 i_127 (.ZN (n_63), .A (p_1[13]));
INV_X1 i_126 (.ZN (n_62), .A (p_1[11]));
OR3_X1 i_125 (.ZN (n_61), .A1 (p_1[2]), .A2 (p_1[1]), .A3 (p_1[0]));
OR2_X1 i_124 (.ZN (n_60), .A1 (n_61), .A2 (p_1[3]));
OR2_X1 i_123 (.ZN (n_59), .A1 (n_60), .A2 (p_1[4]));
OR3_X1 i_122 (.ZN (n_58), .A1 (n_59), .A2 (p_1[5]), .A3 (p_1[6]));
OR2_X1 i_121 (.ZN (n_57), .A1 (n_58), .A2 (p_1[7]));
OR3_X1 i_120 (.ZN (n_56), .A1 (n_57), .A2 (p_1[8]), .A3 (p_1[9]));
NOR2_X1 i_119 (.ZN (n_55), .A1 (n_56), .A2 (p_1[10]));
NAND2_X1 i_118 (.ZN (n_54), .A1 (n_55), .A2 (n_62));
NOR2_X1 i_117 (.ZN (n_53), .A1 (n_54), .A2 (p_1[12]));
NAND2_X1 i_116 (.ZN (n_52), .A1 (n_53), .A2 (n_63));
OR3_X1 i_115 (.ZN (n_51), .A1 (n_52), .A2 (p_1[14]), .A3 (p_1[15]));
OR2_X1 i_114 (.ZN (n_50), .A1 (n_51), .A2 (p_1[16]));
OR2_X1 i_113 (.ZN (n_49), .A1 (n_50), .A2 (p_1[17]));
NOR2_X1 i_112 (.ZN (n_48), .A1 (n_49), .A2 (p_1[18]));
NOR3_X1 i_111 (.ZN (n_47), .A1 (n_49), .A2 (p_1[18]), .A3 (p_1[19]));
NOR4_X1 i_110 (.ZN (n_46), .A1 (n_49), .A2 (p_1[18]), .A3 (p_1[19]), .A4 (p_1[20]));
NAND2_X1 i_109 (.ZN (n_45), .A1 (n_46), .A2 (n_64));
OR2_X1 i_108 (.ZN (n_44), .A1 (n_45), .A2 (p_1[22]));
NOR2_X1 i_107 (.ZN (n_43), .A1 (n_44), .A2 (p_1[23]));
NOR3_X1 i_106 (.ZN (n_42), .A1 (n_44), .A2 (p_1[23]), .A3 (p_1[24]));
NOR4_X1 i_105 (.ZN (n_41), .A1 (n_44), .A2 (p_1[23]), .A3 (p_1[24]), .A4 (p_1[25]));
NAND2_X1 i_104 (.ZN (n_40), .A1 (n_41), .A2 (n_65));
OR2_X1 i_103 (.ZN (n_39), .A1 (n_40), .A2 (p_1[27]));
NOR2_X1 i_102 (.ZN (n_38), .A1 (n_39), .A2 (p_1[28]));
NOR3_X1 i_101 (.ZN (n_37), .A1 (n_39), .A2 (p_1[28]), .A3 (p_1[29]));
NOR4_X1 i_100 (.ZN (n_36), .A1 (n_39), .A2 (p_1[28]), .A3 (p_1[29]), .A4 (p_1[30]));
NAND2_X1 i_99 (.ZN (n_35), .A1 (n_36), .A2 (n_66));
OR2_X1 i_98 (.ZN (n_34), .A1 (n_35), .A2 (p_1[32]));
NOR2_X1 i_97 (.ZN (n_33), .A1 (n_34), .A2 (p_1[33]));
NOR3_X1 i_96 (.ZN (n_32), .A1 (n_34), .A2 (p_1[33]), .A3 (p_1[34]));
NOR4_X1 i_95 (.ZN (n_31), .A1 (n_34), .A2 (p_1[33]), .A3 (p_1[34]), .A4 (p_1[35]));
NAND2_X1 i_94 (.ZN (n_30), .A1 (n_31), .A2 (n_67));
OR2_X1 i_93 (.ZN (n_29), .A1 (n_30), .A2 (p_1[37]));
NOR2_X1 i_92 (.ZN (n_28), .A1 (n_29), .A2 (p_1[38]));
NOR3_X1 i_91 (.ZN (n_27), .A1 (n_29), .A2 (p_1[38]), .A3 (p_1[39]));
NAND2_X1 i_90 (.ZN (n_26), .A1 (n_27), .A2 (n_68));
NOR2_X1 i_89 (.ZN (n_25), .A1 (n_26), .A2 (p_1[41]));
NAND2_X1 i_88 (.ZN (n_24), .A1 (n_25), .A2 (n_69));
OR3_X1 i_87 (.ZN (n_23), .A1 (n_24), .A2 (p_1[43]), .A3 (p_1[44]));
OR2_X1 i_86 (.ZN (n_22), .A1 (n_23), .A2 (p_1[45]));
OR2_X1 i_85 (.ZN (n_21), .A1 (n_22), .A2 (p_1[46]));
OR2_X1 i_84 (.ZN (n_20), .A1 (n_21), .A2 (p_1[47]));
NOR2_X1 i_83 (.ZN (n_19), .A1 (n_20), .A2 (p_1[48]));
NOR3_X1 i_82 (.ZN (n_18), .A1 (n_20), .A2 (p_1[48]), .A3 (p_1[49]));
NOR4_X1 i_81 (.ZN (n_17), .A1 (n_20), .A2 (p_1[48]), .A3 (p_1[49]), .A4 (p_1[50]));
NAND2_X1 i_80 (.ZN (n_16), .A1 (n_17), .A2 (n_70));
NOR2_X1 i_79 (.ZN (n_15), .A1 (n_16), .A2 (p_1[52]));
NOR3_X1 i_78 (.ZN (n_14), .A1 (n_16), .A2 (p_1[52]), .A3 (p_1[53]));
NOR4_X1 i_77 (.ZN (n_13), .A1 (n_16), .A2 (p_1[52]), .A3 (p_1[53]), .A4 (p_1[54]));
NAND2_X1 i_76 (.ZN (n_12), .A1 (n_13), .A2 (n_71));
OR3_X1 i_75 (.ZN (n_11), .A1 (n_12), .A2 (p_1[56]), .A3 (p_1[57]));
NOR2_X1 i_74 (.ZN (n_10), .A1 (n_11), .A2 (p_1[58]));
NOR3_X1 i_73 (.ZN (n_9), .A1 (n_11), .A2 (p_1[58]), .A3 (p_1[59]));
NAND2_X1 i_72 (.ZN (n_8), .A1 (n_9), .A2 (n_72));
NOR2_X1 i_71 (.ZN (n_7), .A1 (n_8), .A2 (p_1[61]));
NOR3_X1 i_70 (.ZN (n_6), .A1 (n_8), .A2 (p_1[61]), .A3 (p_1[62]));
NAND2_X1 i_69 (.ZN (p_0[64]), .A1 (n_6), .A2 (n_73));
XNOR2_X1 i_68 (.ZN (p_0[63]), .A (p_1[63]), .B (n_6));
XNOR2_X1 i_67 (.ZN (p_0[62]), .A (p_1[62]), .B (n_7));
XOR2_X1 i_66 (.Z (p_0[61]), .A (p_1[61]), .B (n_8));
XNOR2_X1 i_65 (.ZN (p_0[60]), .A (p_1[60]), .B (n_9));
XNOR2_X1 i_64 (.ZN (p_0[59]), .A (p_1[59]), .B (n_10));
XOR2_X1 i_63 (.Z (p_0[58]), .A (p_1[58]), .B (n_11));
OAI21_X1 i_62 (.ZN (n_5), .A (p_1[57]), .B1 (n_12), .B2 (p_1[56]));
AND2_X1 i_61 (.ZN (p_0[57]), .A1 (n_11), .A2 (n_5));
XOR2_X1 i_60 (.Z (p_0[56]), .A (p_1[56]), .B (n_12));
XNOR2_X1 i_59 (.ZN (p_0[55]), .A (p_1[55]), .B (n_13));
XNOR2_X1 i_58 (.ZN (p_0[54]), .A (p_1[54]), .B (n_14));
XNOR2_X1 i_57 (.ZN (p_0[53]), .A (p_1[53]), .B (n_15));
XOR2_X1 i_56 (.Z (p_0[52]), .A (p_1[52]), .B (n_16));
XNOR2_X1 i_55 (.ZN (p_0[51]), .A (p_1[51]), .B (n_17));
XNOR2_X1 i_54 (.ZN (p_0[50]), .A (p_1[50]), .B (n_18));
XNOR2_X1 i_53 (.ZN (p_0[49]), .A (p_1[49]), .B (n_19));
XOR2_X1 i_52 (.Z (p_0[48]), .A (p_1[48]), .B (n_20));
XOR2_X1 i_51 (.Z (p_0[47]), .A (p_1[47]), .B (n_21));
XOR2_X1 i_50 (.Z (p_0[46]), .A (p_1[46]), .B (n_22));
XOR2_X1 i_49 (.Z (p_0[45]), .A (p_1[45]), .B (n_23));
OAI21_X1 i_48 (.ZN (n_4), .A (p_1[44]), .B1 (n_24), .B2 (p_1[43]));
AND2_X1 i_47 (.ZN (p_0[44]), .A1 (n_23), .A2 (n_4));
XOR2_X1 i_46 (.Z (p_0[43]), .A (p_1[43]), .B (n_24));
XNOR2_X1 i_45 (.ZN (p_0[42]), .A (p_1[42]), .B (n_25));
XOR2_X1 i_44 (.Z (p_0[41]), .A (p_1[41]), .B (n_26));
XNOR2_X1 i_43 (.ZN (p_0[40]), .A (p_1[40]), .B (n_27));
XNOR2_X1 i_42 (.ZN (p_0[39]), .A (p_1[39]), .B (n_28));
XOR2_X1 i_41 (.Z (p_0[38]), .A (p_1[38]), .B (n_29));
XOR2_X1 i_40 (.Z (p_0[37]), .A (p_1[37]), .B (n_30));
XNOR2_X1 i_39 (.ZN (p_0[36]), .A (p_1[36]), .B (n_31));
XNOR2_X1 i_38 (.ZN (p_0[35]), .A (p_1[35]), .B (n_32));
XNOR2_X1 i_37 (.ZN (p_0[34]), .A (p_1[34]), .B (n_33));
XOR2_X1 i_36 (.Z (p_0[33]), .A (p_1[33]), .B (n_34));
XOR2_X1 i_35 (.Z (p_0[32]), .A (p_1[32]), .B (n_35));
XNOR2_X1 i_34 (.ZN (p_0[31]), .A (p_1[31]), .B (n_36));
XNOR2_X1 i_33 (.ZN (p_0[30]), .A (p_1[30]), .B (n_37));
XNOR2_X1 i_32 (.ZN (p_0[29]), .A (p_1[29]), .B (n_38));
XOR2_X1 i_31 (.Z (p_0[28]), .A (p_1[28]), .B (n_39));
XOR2_X1 i_30 (.Z (p_0[27]), .A (p_1[27]), .B (n_40));
XNOR2_X1 i_29 (.ZN (p_0[26]), .A (p_1[26]), .B (n_41));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (p_1[25]), .B (n_42));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (p_1[24]), .B (n_43));
XOR2_X1 i_26 (.Z (p_0[23]), .A (p_1[23]), .B (n_44));
XOR2_X1 i_25 (.Z (p_0[22]), .A (p_1[22]), .B (n_45));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (p_1[21]), .B (n_46));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (p_1[20]), .B (n_47));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (p_1[19]), .B (n_48));
XOR2_X1 i_21 (.Z (p_0[18]), .A (p_1[18]), .B (n_49));
XOR2_X1 i_20 (.Z (p_0[17]), .A (p_1[17]), .B (n_50));
XOR2_X1 i_19 (.Z (p_0[16]), .A (p_1[16]), .B (n_51));
OAI21_X1 i_18 (.ZN (n_3), .A (p_1[15]), .B1 (n_52), .B2 (p_1[14]));
AND2_X1 i_17 (.ZN (p_0[15]), .A1 (n_51), .A2 (n_3));
XOR2_X1 i_16 (.Z (p_0[14]), .A (p_1[14]), .B (n_52));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (p_1[13]), .B (n_53));
XOR2_X1 i_14 (.Z (p_0[12]), .A (p_1[12]), .B (n_54));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (p_1[11]), .B (n_55));
XOR2_X1 i_12 (.Z (p_0[10]), .A (p_1[10]), .B (n_56));
OAI21_X1 i_11 (.ZN (n_2), .A (p_1[9]), .B1 (n_57), .B2 (p_1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_56), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (p_1[8]), .B (n_57));
XOR2_X1 i_8 (.Z (p_0[7]), .A (p_1[7]), .B (n_58));
OAI21_X1 i_7 (.ZN (n_1), .A (p_1[6]), .B1 (n_59), .B2 (p_1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_58), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (p_1[5]), .B (n_59));
XOR2_X1 i_4 (.Z (p_0[4]), .A (p_1[4]), .B (n_60));
XOR2_X1 i_3 (.Z (p_0[3]), .A (p_1[3]), .B (n_61));
OAI21_X1 i_2 (.ZN (n_0), .A (p_1[2]), .B1 (p_1[1]), .B2 (p_1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_61), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (p_1[1]), .B (p_1[0]));

endmodule //datapath__0_11

module datapath__0_9 (m, p_0, p_1);

output [32:0] p_1;
input [31:0] m;
input [31:0] p_0;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;


FA_X1 i_31 (.CO (p_1[32]), .S (p_1[31]), .A (m[31]), .B (p_0[31]), .CI (n_30));
FA_X1 i_30 (.CO (n_30), .S (p_1[30]), .A (m[30]), .B (p_0[30]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_1[29]), .A (m[29]), .B (p_0[29]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_1[28]), .A (m[28]), .B (p_0[28]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_1[27]), .A (m[27]), .B (p_0[27]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_1[26]), .A (m[26]), .B (p_0[26]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_1[25]), .A (m[25]), .B (p_0[25]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_1[24]), .A (m[24]), .B (p_0[24]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_1[23]), .A (m[23]), .B (p_0[23]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_1[22]), .A (m[22]), .B (p_0[22]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_1[21]), .A (m[21]), .B (p_0[21]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_1[20]), .A (m[20]), .B (p_0[20]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_1[19]), .A (m[19]), .B (p_0[19]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_1[18]), .A (m[18]), .B (p_0[18]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_1[17]), .A (m[17]), .B (p_0[17]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_1[16]), .A (m[16]), .B (p_0[16]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_1[15]), .A (m[15]), .B (p_0[15]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_1[14]), .A (m[14]), .B (p_0[14]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_1[13]), .A (m[13]), .B (p_0[13]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_1[12]), .A (m[12]), .B (p_0[12]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_1[11]), .A (m[11]), .B (p_0[11]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_1[10]), .A (m[10]), .B (p_0[10]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_1[9]), .A (m[9]), .B (p_0[9]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_1[8]), .A (m[8]), .B (p_0[8]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_1[7]), .A (m[7]), .B (p_0[7]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_1[6]), .A (m[6]), .B (p_0[6]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_1[5]), .A (m[5]), .B (p_0[5]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_1[4]), .A (m[4]), .B (p_0[4]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_1[3]), .A (m[3]), .B (p_0[3]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_1[2]), .A (m[2]), .B (p_0[2]), .CI (n_1));
FA_X1 i_1 (.CO (n_1), .S (p_1[1]), .A (m[1]), .B (p_0[1]), .CI (n_0));
HA_X1 i_0 (.CO (n_0), .S (p_1[0]), .A (m[0]), .B (p_0[0]));

endmodule //datapath__0_9

module datapath__0_2 (p_0, in1);

output [31:0] p_0;
input [31:0] in1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (in1[25]));
INV_X1 i_63 (.ZN (n_32), .A (in1[21]));
INV_X1 i_62 (.ZN (n_31), .A (in1[14]));
INV_X1 i_61 (.ZN (n_30), .A (in1[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (in1[2]), .A2 (in1[1]), .A3 (in1[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (in1[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (in1[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (in1[5]), .A3 (in1[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (in1[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (in1[8]), .A3 (in1[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (in1[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (in1[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (in1[12]), .A3 (in1[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (in1[15]), .A3 (in1[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (in1[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (in1[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (in1[18]), .A3 (in1[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (in1[18]), .A3 (in1[19]), .A4 (in1[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (in1[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (in1[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (in1[23]), .A3 (in1[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (in1[26]), .A3 (in1[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (in1[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (in1[28]), .A3 (in1[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (in1[28]), .A3 (in1[29]), .A4 (in1[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (in1[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (in1[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (in1[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (in1[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (in1[27]), .B1 (n_9), .B2 (in1[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (in1[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (in1[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (in1[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (in1[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (in1[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (in1[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (in1[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (in1[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (in1[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (in1[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (in1[16]), .B1 (n_19), .B2 (in1[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (in1[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (in1[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (in1[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (in1[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (in1[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (in1[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (in1[9]), .B1 (n_25), .B2 (in1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (in1[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (in1[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (in1[6]), .B1 (n_27), .B2 (in1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (in1[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (in1[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (in1[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (in1[2]), .B1 (in1[1]), .B2 (in1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (in1[1]), .B (in1[0]));

endmodule //datapath__0_2

module datapath (p_0, in2);

output [31:0] p_0;
input [31:0] in2;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (in2[25]));
INV_X1 i_63 (.ZN (n_32), .A (in2[21]));
INV_X1 i_62 (.ZN (n_31), .A (in2[14]));
INV_X1 i_61 (.ZN (n_30), .A (in2[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (in2[2]), .A2 (in2[1]), .A3 (in2[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (in2[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (in2[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (in2[5]), .A3 (in2[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (in2[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (in2[8]), .A3 (in2[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (in2[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (in2[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (in2[12]), .A3 (in2[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (in2[15]), .A3 (in2[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (in2[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (in2[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (in2[18]), .A3 (in2[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (in2[18]), .A3 (in2[19]), .A4 (in2[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (in2[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (in2[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (in2[23]), .A3 (in2[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (in2[26]), .A3 (in2[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (in2[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (in2[28]), .A3 (in2[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (in2[28]), .A3 (in2[29]), .A4 (in2[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (in2[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (in2[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (in2[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (in2[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (in2[27]), .B1 (n_9), .B2 (in2[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (in2[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (in2[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (in2[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (in2[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (in2[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (in2[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (in2[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (in2[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (in2[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (in2[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (in2[16]), .B1 (n_19), .B2 (in2[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (in2[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (in2[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (in2[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (in2[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (in2[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (in2[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (in2[9]), .B1 (n_25), .B2 (in2[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (in2[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (in2[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (in2[6]), .B1 (n_27), .B2 (in2[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (in2[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (in2[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (in2[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (in2[2]), .B1 (in2[1]), .B2 (in2[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (in2[1]), .B (in2[0]));

endmodule //datapath

module sequentialmultiplier (clk_CTS_0_PP_1, clk_CTS_0_PP_0, clk_CTS_0_PP_15, CTSclk_CTS_0_PP_15PP_0, 
    in1, in2, clk, reset, en, result, enableOutput);

output enableOutput;
output [63:0] result;
output clk_CTS_0_PP_1;
input clk;
input en;
input [31:0] in1;
input [31:0] in2;
input reset;
input clk_CTS_0_PP_0;
input clk_CTS_0_PP_15;
input CTSclk_CTS_0_PP_15PP_0;
wire CTS_n_tid0_179;
wire \counter[5] ;
wire \counter[4] ;
wire \counter[3] ;
wire \counter[2] ;
wire \counter[1] ;
wire \counter[0] ;
wire resetReg;
wire \res[64] ;
wire \res[63] ;
wire \res[62] ;
wire \res[61] ;
wire \res[60] ;
wire \res[59] ;
wire \res[58] ;
wire \res[57] ;
wire \res[56] ;
wire \res[55] ;
wire \res[54] ;
wire \res[53] ;
wire \res[52] ;
wire \res[51] ;
wire \res[50] ;
wire \res[49] ;
wire \res[48] ;
wire \res[47] ;
wire \res[46] ;
wire \res[45] ;
wire \res[44] ;
wire \res[43] ;
wire \res[42] ;
wire \res[41] ;
wire \res[40] ;
wire \res[39] ;
wire \res[38] ;
wire \res[37] ;
wire \res[36] ;
wire \res[35] ;
wire \res[34] ;
wire \res[33] ;
wire \res[32] ;
wire \res[31] ;
wire \res[30] ;
wire \res[29] ;
wire \res[28] ;
wire \res[27] ;
wire \res[26] ;
wire \res[25] ;
wire \res[24] ;
wire \res[23] ;
wire \res[22] ;
wire \res[21] ;
wire \res[20] ;
wire \res[19] ;
wire \res[18] ;
wire \res[17] ;
wire \res[16] ;
wire \res[15] ;
wire \res[14] ;
wire \res[13] ;
wire \res[12] ;
wire \res[11] ;
wire \res[10] ;
wire \res[9] ;
wire \res[8] ;
wire \res[7] ;
wire \res[6] ;
wire \res[5] ;
wire \res[4] ;
wire \res[3] ;
wire \res[2] ;
wire \res[1] ;
wire \res[0] ;
wire n_1_3;
wire n_1_0;
wire n_1_4;
wire n_1_1;
wire n_1_5;
wire n_1_2;
wire n_1_6;
wire n_1_7;
wire n_1_8;
wire n_1_9;
wire n_1_10;
wire n_1_11;
wire n_1_12;
wire n_1_13;
wire n_1_14;
wire n_1_15;
wire n_1_16;
wire n_1_17;
wire n_1_18;
wire n_1_19;
wire n_1_20;
wire n_1_21;
wire n_1_22;
wire n_1_23;
wire n_1_24;
wire n_1_25;
wire n_1_26;
wire n_1_27;
wire n_1_28;
wire n_1_29;
wire n_1_30;
wire n_1_31;
wire n_1_32;
wire n_1_33;
wire n_1_34;
wire n_1_35;
wire n_1_36;
wire n_1_37;
wire n_1_38;
wire n_1_39;
wire n_1_40;
wire n_1_41;
wire n_1_42;
wire n_1_43;
wire n_1_44;
wire n_1_45;
wire n_1_46;
wire n_1_47;
wire n_1_48;
wire n_1_49;
wire n_1_50;
wire n_1_51;
wire n_1_52;
wire n_1_53;
wire n_1_54;
wire n_1_55;
wire n_1_56;
wire n_1_57;
wire n_1_58;
wire n_1_59;
wire n_1_60;
wire n_1_61;
wire n_1_62;
wire n_1_63;
wire n_1_64;
wire n_1_65;
wire n_1_66;
wire n_1_67;
wire n_1_68;
wire n_1_69;
wire n_1_70;
wire n_1_71;
wire n_1_72;
wire n_1_73;
wire n_1_74;
wire n_1_75;
wire n_1_76;
wire n_1_77;
wire n_1_78;
wire n_1_79;
wire n_1_80;
wire n_1_81;
wire n_1_83;
wire n_1_84;
wire n_1_85;
wire n_1_86;
wire n_1_87;
wire n_1_88;
wire n_1_89;
wire n_1_90;
wire n_1_91;
wire n_1_92;
wire n_1_93;
wire n_1_94;
wire n_1_95;
wire n_1_96;
wire n_1_97;
wire n_1_98;
wire n_1_99;
wire n_1_100;
wire n_1_101;
wire n_1_102;
wire n_1_103;
wire n_1_104;
wire n_1_105;
wire n_1_106;
wire n_1_107;
wire n_1_108;
wire n_1_109;
wire n_1_110;
wire n_1_111;
wire n_1_112;
wire n_1_113;
wire n_1_114;
wire n_1_115;
wire n_1_116;
wire n_1_117;
wire n_1_118;
wire n_1_119;
wire n_1_120;
wire n_1_121;
wire n_1_122;
wire n_1_123;
wire n_1_124;
wire n_1_125;
wire n_1_126;
wire n_1_127;
wire n_1_128;
wire n_1_129;
wire n_1_130;
wire n_1_131;
wire n_1_132;
wire n_1_133;
wire n_1_134;
wire n_1_135;
wire n_1_136;
wire n_1_137;
wire n_1_138;
wire n_1_139;
wire n_1_140;
wire n_1_141;
wire n_1_142;
wire n_1_143;
wire n_1_144;
wire n_1_145;
wire n_1_146;
wire n_1_147;
wire n_1_148;
wire n_1_149;
wire n_1_150;
wire n_1_151;
wire n_1_152;
wire n_1_153;
wire n_1_154;
wire n_1_155;
wire n_1_156;
wire n_1_157;
wire n_1_158;
wire n_1_159;
wire n_1_160;
wire n_1_161;
wire n_1_162;
wire n_1_163;
wire n_1_164;
wire n_1_165;
wire n_1_166;
wire n_1_167;
wire n_1_168;
wire n_1_169;
wire n_1_170;
wire n_1_171;
wire n_1_184;
wire \m[31] ;
wire \m[30] ;
wire \m[29] ;
wire \m[28] ;
wire \m[27] ;
wire \m[26] ;
wire \m[25] ;
wire \m[24] ;
wire \m[23] ;
wire \m[22] ;
wire \m[21] ;
wire \m[20] ;
wire \m[19] ;
wire \m[18] ;
wire \m[17] ;
wire \m[16] ;
wire \m[15] ;
wire \m[14] ;
wire \m[13] ;
wire \m[12] ;
wire \m[11] ;
wire \m[10] ;
wire \m[9] ;
wire \m[8] ;
wire \m[7] ;
wire \m[6] ;
wire \m[5] ;
wire \m[4] ;
wire \m[3] ;
wire \m[2] ;
wire \m[1] ;
wire hfn_ipo_n22;
wire n_1_188;
wire n_1_82;
wire n_1_172;
wire n_1_173;
wire n_1_174;
wire n_1_175;
wire n_1_176;
wire n_1_177;
wire n_1_178;
wire n_1_179;
wire n_1_180;
wire n_1_181;
wire n_1_182;
wire n_1_183;
wire n_1_185;
wire n_1_186;
wire n_1_187;
wire n_1_189;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire uc_0;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire uc_1;
wire n_334;
wire n_97;
wire n_96;
wire n_95;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_161;
wire n_160;
wire n_159;
wire n_158;
wire n_157;
wire n_156;
wire n_155;
wire n_154;
wire n_153;
wire n_152;
wire n_151;
wire n_150;
wire n_149;
wire n_148;
wire n_147;
wire n_146;
wire n_145;
wire n_144;
wire n_143;
wire n_142;
wire n_141;
wire n_140;
wire n_139;
wire n_138;
wire n_137;
wire n_136;
wire n_135;
wire n_134;
wire n_133;
wire n_132;
wire n_131;
wire n_130;
wire n_129;
wire n_128;
wire n_127;
wire n_126;
wire n_125;
wire n_124;
wire n_123;
wire n_122;
wire n_121;
wire n_120;
wire n_119;
wire n_118;
wire n_117;
wire n_116;
wire n_115;
wire n_114;
wire n_113;
wire n_112;
wire n_111;
wire n_110;
wire n_109;
wire n_108;
wire n_107;
wire n_106;
wire n_105;
wire n_104;
wire n_103;
wire n_102;
wire n_101;
wire n_100;
wire n_99;
wire n_98;
wire uc_2;
wire n_331;
wire n_330;
wire n_329;
wire n_328;
wire n_327;
wire n_326;
wire n_325;
wire n_324;
wire n_323;
wire n_322;
wire n_321;
wire n_320;
wire n_319;
wire n_318;
wire n_317;
wire n_316;
wire n_315;
wire n_314;
wire n_313;
wire n_312;
wire n_311;
wire n_310;
wire n_309;
wire n_308;
wire n_307;
wire n_306;
wire n_305;
wire n_304;
wire n_303;
wire n_302;
wire n_301;
wire n_300;
wire n_299;
wire n_333;
wire CTS_n_tid0_91;
wire n_227;
wire n_226;
wire n_225;
wire n_224;
wire n_223;
wire n_222;
wire n_221;
wire n_220;
wire n_219;
wire n_218;
wire n_217;
wire n_216;
wire n_215;
wire n_214;
wire n_213;
wire n_212;
wire n_211;
wire n_210;
wire n_209;
wire n_208;
wire n_207;
wire n_206;
wire n_205;
wire n_204;
wire n_203;
wire n_202;
wire n_201;
wire n_200;
wire n_199;
wire n_198;
wire n_197;
wire n_196;
wire n_195;
wire n_194;
wire n_193;
wire n_192;
wire n_191;
wire n_190;
wire n_189;
wire n_188;
wire n_187;
wire n_186;
wire n_185;
wire n_184;
wire n_183;
wire n_182;
wire n_181;
wire n_180;
wire n_179;
wire n_178;
wire n_177;
wire n_176;
wire n_175;
wire n_174;
wire n_173;
wire n_172;
wire n_171;
wire n_170;
wire n_169;
wire n_168;
wire n_167;
wire n_166;
wire n_165;
wire n_164;
wire n_1;
wire n_233;
wire n_232;
wire n_231;
wire n_230;
wire n_229;
wire n_228;
wire n_162;
wire n_163;
wire n_335;
wire n_332;
wire CTS_n_tid1_32;
wire n_298;
wire n_297;
wire n_296;
wire n_295;
wire n_294;
wire n_293;
wire n_292;
wire n_291;
wire n_290;
wire n_289;
wire n_288;
wire n_287;
wire n_286;
wire n_285;
wire n_284;
wire n_283;
wire n_282;
wire n_281;
wire n_280;
wire n_279;
wire n_278;
wire n_277;
wire n_276;
wire n_275;
wire n_274;
wire n_273;
wire n_272;
wire n_271;
wire n_270;
wire n_269;
wire n_268;
wire n_267;
wire n_266;
wire n_265;
wire n_264;
wire n_263;
wire n_262;
wire n_261;
wire n_260;
wire n_259;
wire n_258;
wire n_257;
wire n_256;
wire n_255;
wire n_254;
wire n_253;
wire n_252;
wire n_251;
wire n_250;
wire n_249;
wire n_248;
wire n_247;
wire n_246;
wire n_245;
wire n_244;
wire n_243;
wire n_242;
wire n_241;
wire n_240;
wire n_239;
wire n_238;
wire n_237;
wire n_236;
wire n_235;
wire n_234;
wire hfn_ipo_n23;
wire hfn_ipo_n24;
wire hfn_ipo_n25;
wire hfn_ipo_n27;
wire hfn_ipo_n28;
wire drc_ipo_n29;
wire drc_ipo_n30;
wire hfn_ipo_n26;
wire hfn_ipo_n21;
wire CTS_n_tid1_33;
wire CTS_n_tid0_92;
wire CTS_n_tid1_82;


INV_X1 i_1_389 (.ZN (n_1_189), .A (\counter[5] ));
INV_X1 i_1_388 (.ZN (n_1_187), .A (n_1_6));
NOR4_X1 i_1_387 (.ZN (n_1_186), .A1 (\counter[4] ), .A2 (\counter[3] ), .A3 (\counter[2] ), .A4 (\counter[1] ));
INV_X1 i_1_386 (.ZN (n_1_185), .A (n_1_186));
NOR2_X1 i_1_373 (.ZN (n_1_183), .A1 (\counter[0] ), .A2 (n_1_185));
OAI21_X1 i_1_372 (.ZN (n_1_182), .A (n_1_183), .B1 (n_1_189), .B2 (\counter[4] ));
INV_X1 i_1_354 (.ZN (n_1_181), .A (n_1_182));
NOR3_X1 i_1_353 (.ZN (n_1_180), .A1 (reset), .A2 (resetReg), .A3 (n_1_181));
INV_X1 i_1_352 (.ZN (n_1_179), .A (n_1_180));
XOR2_X1 i_1_351 (.Z (n_1_178), .A (\counter[5] ), .B (n_1_7));
NOR3_X1 i_1_350 (.ZN (n_1_177), .A1 (n_1_5), .A2 (n_1_4), .A3 (n_1_3));
NAND4_X1 i_1_349 (.ZN (n_1_176), .A1 (\counter[0] ), .A2 (n_1_187), .A3 (n_1_177), .A4 (n_1_178));
XNOR2_X1 i_1_348 (.ZN (n_1_175), .A (in2[31]), .B (in1[31]));
NOR2_X1 i_1_347 (.ZN (n_1_174), .A1 (n_1_176), .A2 (n_1_175));
NOR2_X1 i_1_346 (.ZN (n_1_173), .A1 (n_1_179), .A2 (n_1_174));
AND2_X1 i_1_345 (.ZN (n_1_172), .A1 (n_1_180), .A2 (n_1_174));
AOI22_X1 i_1_331 (.ZN (n_1_82), .A1 (\res[5] ), .A2 (hfn_ipo_n28), .B1 (n_101), .B2 (hfn_ipo_n26));
INV_X1 i_1_330 (.ZN (n_1_188), .A (en));
AND2_X1 i_1_385 (.ZN (\m[31] ), .A1 (in1[31]), .A2 (n_64));
MUX2_X1 i_1_384 (.Z (\m[30] ), .A (in1[30]), .B (n_63), .S (in1[31]));
MUX2_X1 i_1_383 (.Z (\m[29] ), .A (in1[29]), .B (n_62), .S (in1[31]));
MUX2_X1 i_1_382 (.Z (\m[28] ), .A (in1[28]), .B (n_61), .S (in1[31]));
MUX2_X1 i_1_381 (.Z (\m[27] ), .A (in1[27]), .B (n_60), .S (in1[31]));
MUX2_X1 i_1_380 (.Z (\m[26] ), .A (in1[26]), .B (n_59), .S (in1[31]));
MUX2_X1 i_1_379 (.Z (\m[25] ), .A (in1[25]), .B (n_58), .S (in1[31]));
MUX2_X1 i_1_378 (.Z (\m[24] ), .A (in1[24]), .B (n_57), .S (in1[31]));
MUX2_X1 i_1_377 (.Z (\m[23] ), .A (in1[23]), .B (n_56), .S (in1[31]));
MUX2_X1 i_1_376 (.Z (\m[22] ), .A (in1[22]), .B (n_55), .S (in1[31]));
MUX2_X1 i_1_375 (.Z (\m[21] ), .A (in1[21]), .B (n_54), .S (in1[31]));
MUX2_X1 i_1_374 (.Z (\m[20] ), .A (in1[20]), .B (n_53), .S (in1[31]));
MUX2_X1 i_1_329 (.Z (\m[19] ), .A (in1[19]), .B (n_52), .S (in1[31]));
MUX2_X1 i_1_328 (.Z (\m[18] ), .A (in1[18]), .B (n_51), .S (in1[31]));
MUX2_X1 i_1_371 (.Z (\m[17] ), .A (in1[17]), .B (n_50), .S (in1[31]));
MUX2_X1 i_1_370 (.Z (\m[16] ), .A (in1[16]), .B (n_49), .S (in1[31]));
MUX2_X1 i_1_369 (.Z (\m[15] ), .A (in1[15]), .B (n_48), .S (in1[31]));
MUX2_X1 i_1_368 (.Z (\m[14] ), .A (in1[14]), .B (n_47), .S (in1[31]));
MUX2_X1 i_1_367 (.Z (\m[13] ), .A (in1[13]), .B (n_46), .S (in1[31]));
MUX2_X1 i_1_366 (.Z (\m[12] ), .A (in1[12]), .B (n_45), .S (in1[31]));
MUX2_X1 i_1_365 (.Z (\m[11] ), .A (in1[11]), .B (n_44), .S (in1[31]));
MUX2_X1 i_1_364 (.Z (\m[10] ), .A (in1[10]), .B (n_43), .S (in1[31]));
MUX2_X1 i_1_363 (.Z (\m[9] ), .A (in1[9]), .B (n_42), .S (in1[31]));
MUX2_X1 i_1_362 (.Z (\m[8] ), .A (in1[8]), .B (n_41), .S (in1[31]));
MUX2_X1 i_1_361 (.Z (\m[7] ), .A (in1[7]), .B (n_40), .S (in1[31]));
MUX2_X1 i_1_360 (.Z (\m[6] ), .A (in1[6]), .B (n_39), .S (in1[31]));
MUX2_X1 i_1_359 (.Z (\m[5] ), .A (in1[5]), .B (n_38), .S (in1[31]));
MUX2_X1 i_1_358 (.Z (\m[4] ), .A (in1[4]), .B (n_37), .S (in1[31]));
MUX2_X1 i_1_357 (.Z (\m[3] ), .A (in1[3]), .B (n_36), .S (in1[31]));
MUX2_X1 i_1_356 (.Z (\m[2] ), .A (in1[2]), .B (n_35), .S (in1[31]));
MUX2_X1 i_1_355 (.Z (\m[1] ), .A (in1[1]), .B (n_34), .S (in1[31]));
OAI21_X1 i_1_311 (.ZN (n_1_184), .A (en), .B1 (reset), .B2 (resetReg));
INV_X1 i_1_310 (.ZN (n_335), .A (n_1_184));
AOI21_X1 i_1_309 (.ZN (n_334), .A (n_335), .B1 (n_1_176), .B2 (en));
NAND2_X1 i_1_308 (.ZN (n_333), .A1 (n_1_184), .A2 (n_1_176));
NOR3_X1 i_1_307 (.ZN (n_332), .A1 (n_1_188), .A2 (reset), .A3 (resetReg));
MUX2_X1 i_1_344 (.Z (n_331), .A (\res[64] ), .B (n_97), .S (drc_ipo_n30));
MUX2_X1 i_1_343 (.Z (n_330), .A (\res[63] ), .B (n_96), .S (drc_ipo_n30));
MUX2_X1 i_1_342 (.Z (n_329), .A (\res[62] ), .B (n_95), .S (drc_ipo_n30));
MUX2_X1 i_1_341 (.Z (n_328), .A (\res[61] ), .B (n_94), .S (drc_ipo_n30));
MUX2_X1 i_1_340 (.Z (n_327), .A (\res[60] ), .B (n_93), .S (drc_ipo_n30));
MUX2_X1 i_1_339 (.Z (n_326), .A (\res[59] ), .B (n_92), .S (drc_ipo_n30));
MUX2_X1 i_1_338 (.Z (n_325), .A (\res[58] ), .B (n_91), .S (drc_ipo_n30));
MUX2_X1 i_1_337 (.Z (n_324), .A (\res[57] ), .B (n_90), .S (drc_ipo_n30));
MUX2_X1 i_1_336 (.Z (n_323), .A (\res[56] ), .B (n_89), .S (drc_ipo_n30));
MUX2_X1 i_1_335 (.Z (n_322), .A (\res[55] ), .B (n_88), .S (drc_ipo_n30));
MUX2_X1 i_1_334 (.Z (n_321), .A (\res[54] ), .B (n_87), .S (drc_ipo_n30));
MUX2_X1 i_1_333 (.Z (n_320), .A (\res[53] ), .B (n_86), .S (drc_ipo_n30));
MUX2_X1 i_1_332 (.Z (n_319), .A (\res[52] ), .B (n_85), .S (drc_ipo_n30));
MUX2_X1 i_1_306 (.Z (n_318), .A (\res[51] ), .B (n_84), .S (drc_ipo_n30));
MUX2_X1 i_1_304 (.Z (n_317), .A (\res[50] ), .B (n_83), .S (drc_ipo_n30));
MUX2_X1 i_1_303 (.Z (n_316), .A (\res[49] ), .B (n_82), .S (drc_ipo_n30));
MUX2_X1 i_1_300 (.Z (n_315), .A (\res[48] ), .B (n_81), .S (drc_ipo_n30));
MUX2_X1 i_1_327 (.Z (n_314), .A (\res[47] ), .B (n_80), .S (drc_ipo_n30));
MUX2_X1 i_1_326 (.Z (n_313), .A (\res[46] ), .B (n_79), .S (drc_ipo_n30));
MUX2_X1 i_1_325 (.Z (n_312), .A (\res[45] ), .B (n_78), .S (drc_ipo_n30));
MUX2_X1 i_1_324 (.Z (n_311), .A (\res[44] ), .B (n_77), .S (drc_ipo_n30));
MUX2_X1 i_1_323 (.Z (n_310), .A (\res[43] ), .B (n_76), .S (drc_ipo_n30));
MUX2_X1 i_1_322 (.Z (n_309), .A (\res[42] ), .B (n_75), .S (drc_ipo_n30));
MUX2_X1 i_1_321 (.Z (n_308), .A (\res[41] ), .B (n_74), .S (drc_ipo_n30));
MUX2_X1 i_1_320 (.Z (n_307), .A (\res[40] ), .B (n_73), .S (drc_ipo_n30));
MUX2_X1 i_1_319 (.Z (n_306), .A (\res[39] ), .B (n_72), .S (drc_ipo_n30));
MUX2_X1 i_1_318 (.Z (n_305), .A (\res[38] ), .B (n_71), .S (drc_ipo_n30));
MUX2_X1 i_1_317 (.Z (n_304), .A (\res[37] ), .B (n_70), .S (drc_ipo_n30));
MUX2_X1 i_1_316 (.Z (n_303), .A (\res[36] ), .B (n_69), .S (drc_ipo_n30));
MUX2_X1 i_1_315 (.Z (n_302), .A (\res[35] ), .B (n_68), .S (drc_ipo_n30));
MUX2_X1 i_1_314 (.Z (n_301), .A (\res[34] ), .B (n_67), .S (drc_ipo_n30));
MUX2_X1 i_1_313 (.Z (n_300), .A (\res[33] ), .B (n_66), .S (drc_ipo_n30));
MUX2_X1 i_1_312 (.Z (n_299), .A (\res[32] ), .B (n_65), .S (drc_ipo_n30));
AND3_X1 i_1_305 (.ZN (n_298), .A1 (n_161), .A2 (n_1_180), .A3 (n_1_174));
AOI22_X1 i_1_302 (.ZN (n_1_171), .A1 (n_160), .A2 (hfn_ipo_n26), .B1 (hfn_ipo_n28), .B2 (n_331));
INV_X1 i_1_301 (.ZN (n_297), .A (n_1_171));
NOR3_X1 i_1_299 (.ZN (n_1_170), .A1 (n_1_182), .A2 (resetReg), .A3 (reset));
AND2_X2 i_1_274 (.ZN (n_1_169), .A1 (in2[0]), .A2 (n_1_170));
AOI222_X1 i_1_298 (.ZN (n_1_168), .A1 (n_159), .A2 (hfn_ipo_n26), .B1 (n_1_169), .B2 (\m[31] )
    , .C1 (n_330), .C2 (hfn_ipo_n28));
INV_X1 i_1_297 (.ZN (n_296), .A (n_1_168));
AOI222_X1 i_1_296 (.ZN (n_1_167), .A1 (n_1_169), .A2 (\m[30] ), .B1 (n_158), .B2 (hfn_ipo_n26)
    , .C1 (n_329), .C2 (hfn_ipo_n28));
INV_X1 i_1_295 (.ZN (n_295), .A (n_1_167));
AOI222_X1 i_1_294 (.ZN (n_1_166), .A1 (n_1_169), .A2 (\m[29] ), .B1 (n_157), .B2 (hfn_ipo_n26)
    , .C1 (n_328), .C2 (hfn_ipo_n28));
INV_X1 i_1_293 (.ZN (n_294), .A (n_1_166));
AOI222_X1 i_1_292 (.ZN (n_1_165), .A1 (n_1_169), .A2 (\m[28] ), .B1 (n_156), .B2 (hfn_ipo_n26)
    , .C1 (n_327), .C2 (hfn_ipo_n28));
INV_X1 i_1_291 (.ZN (n_293), .A (n_1_165));
AOI222_X1 i_1_290 (.ZN (n_1_164), .A1 (n_1_169), .A2 (\m[27] ), .B1 (n_155), .B2 (hfn_ipo_n26)
    , .C1 (n_326), .C2 (hfn_ipo_n28));
INV_X1 i_1_289 (.ZN (n_292), .A (n_1_164));
AOI222_X1 i_1_288 (.ZN (n_1_163), .A1 (n_1_169), .A2 (\m[26] ), .B1 (n_154), .B2 (hfn_ipo_n26)
    , .C1 (n_325), .C2 (hfn_ipo_n28));
INV_X1 i_1_287 (.ZN (n_291), .A (n_1_163));
AOI222_X1 i_1_286 (.ZN (n_1_162), .A1 (n_1_169), .A2 (\m[25] ), .B1 (n_153), .B2 (hfn_ipo_n26)
    , .C1 (n_324), .C2 (hfn_ipo_n28));
INV_X1 i_1_285 (.ZN (n_290), .A (n_1_162));
AOI222_X1 i_1_284 (.ZN (n_1_161), .A1 (n_1_169), .A2 (\m[24] ), .B1 (n_152), .B2 (hfn_ipo_n26)
    , .C1 (n_323), .C2 (hfn_ipo_n28));
INV_X1 i_1_283 (.ZN (n_289), .A (n_1_161));
AOI222_X1 i_1_282 (.ZN (n_1_160), .A1 (n_1_169), .A2 (\m[23] ), .B1 (n_151), .B2 (hfn_ipo_n26)
    , .C1 (n_322), .C2 (hfn_ipo_n28));
INV_X1 i_1_281 (.ZN (n_288), .A (n_1_160));
AOI222_X1 i_1_280 (.ZN (n_1_159), .A1 (n_1_169), .A2 (\m[22] ), .B1 (n_150), .B2 (hfn_ipo_n26)
    , .C1 (n_321), .C2 (hfn_ipo_n28));
INV_X1 i_1_279 (.ZN (n_287), .A (n_1_159));
AOI222_X1 i_1_278 (.ZN (n_1_158), .A1 (n_1_169), .A2 (\m[21] ), .B1 (n_149), .B2 (hfn_ipo_n26)
    , .C1 (n_320), .C2 (hfn_ipo_n28));
INV_X1 i_1_277 (.ZN (n_286), .A (n_1_158));
AOI222_X1 i_1_276 (.ZN (n_1_157), .A1 (n_1_169), .A2 (\m[20] ), .B1 (n_148), .B2 (hfn_ipo_n26)
    , .C1 (n_319), .C2 (hfn_ipo_n28));
INV_X1 i_1_275 (.ZN (n_285), .A (n_1_157));
AOI222_X1 i_1_273 (.ZN (n_1_156), .A1 (n_1_169), .A2 (\m[19] ), .B1 (n_147), .B2 (hfn_ipo_n26)
    , .C1 (n_318), .C2 (hfn_ipo_n28));
INV_X1 i_1_272 (.ZN (n_284), .A (n_1_156));
AOI222_X1 i_1_233 (.ZN (n_1_155), .A1 (n_1_169), .A2 (\m[18] ), .B1 (n_146), .B2 (hfn_ipo_n26)
    , .C1 (n_317), .C2 (hfn_ipo_n28));
INV_X1 i_1_271 (.ZN (n_283), .A (n_1_155));
AOI222_X1 i_1_270 (.ZN (n_1_154), .A1 (n_1_169), .A2 (\m[17] ), .B1 (n_145), .B2 (hfn_ipo_n26)
    , .C1 (n_316), .C2 (hfn_ipo_n28));
INV_X1 i_1_269 (.ZN (n_282), .A (n_1_154));
AOI222_X1 i_1_268 (.ZN (n_1_153), .A1 (n_1_169), .A2 (\m[16] ), .B1 (n_144), .B2 (hfn_ipo_n26)
    , .C1 (n_315), .C2 (hfn_ipo_n28));
INV_X1 i_1_267 (.ZN (n_281), .A (n_1_153));
AOI222_X1 i_1_266 (.ZN (n_1_152), .A1 (n_1_169), .A2 (\m[15] ), .B1 (n_143), .B2 (hfn_ipo_n26)
    , .C1 (n_314), .C2 (hfn_ipo_n28));
INV_X1 i_1_265 (.ZN (n_280), .A (n_1_152));
AOI222_X1 i_1_264 (.ZN (n_1_151), .A1 (n_1_169), .A2 (\m[14] ), .B1 (n_142), .B2 (hfn_ipo_n26)
    , .C1 (n_313), .C2 (hfn_ipo_n28));
INV_X1 i_1_263 (.ZN (n_279), .A (n_1_151));
AOI222_X1 i_1_262 (.ZN (n_1_150), .A1 (n_1_169), .A2 (\m[13] ), .B1 (n_141), .B2 (hfn_ipo_n26)
    , .C1 (n_312), .C2 (hfn_ipo_n28));
INV_X1 i_1_261 (.ZN (n_278), .A (n_1_150));
AOI222_X1 i_1_260 (.ZN (n_1_149), .A1 (n_1_169), .A2 (\m[12] ), .B1 (n_140), .B2 (hfn_ipo_n26)
    , .C1 (n_311), .C2 (hfn_ipo_n28));
INV_X1 i_1_259 (.ZN (n_277), .A (n_1_149));
AOI222_X1 i_1_258 (.ZN (n_1_148), .A1 (n_1_169), .A2 (\m[11] ), .B1 (n_139), .B2 (hfn_ipo_n26)
    , .C1 (n_310), .C2 (hfn_ipo_n28));
INV_X1 i_1_257 (.ZN (n_276), .A (n_1_148));
AOI222_X1 i_1_256 (.ZN (n_1_147), .A1 (n_1_169), .A2 (\m[10] ), .B1 (n_138), .B2 (hfn_ipo_n26)
    , .C1 (n_309), .C2 (hfn_ipo_n28));
INV_X1 i_1_255 (.ZN (n_275), .A (n_1_147));
AOI222_X1 i_1_254 (.ZN (n_1_146), .A1 (n_1_169), .A2 (\m[9] ), .B1 (n_137), .B2 (hfn_ipo_n26)
    , .C1 (n_308), .C2 (hfn_ipo_n28));
INV_X1 i_1_253 (.ZN (n_274), .A (n_1_146));
AOI222_X1 i_1_252 (.ZN (n_1_145), .A1 (n_1_169), .A2 (\m[8] ), .B1 (n_136), .B2 (hfn_ipo_n25)
    , .C1 (n_307), .C2 (hfn_ipo_n27));
INV_X1 i_1_251 (.ZN (n_273), .A (n_1_145));
AOI222_X1 i_1_250 (.ZN (n_1_144), .A1 (n_1_169), .A2 (\m[7] ), .B1 (n_135), .B2 (hfn_ipo_n25)
    , .C1 (n_306), .C2 (hfn_ipo_n27));
INV_X1 i_1_249 (.ZN (n_272), .A (n_1_144));
AOI222_X1 i_1_248 (.ZN (n_1_143), .A1 (n_1_169), .A2 (\m[6] ), .B1 (n_134), .B2 (hfn_ipo_n25)
    , .C1 (n_305), .C2 (hfn_ipo_n27));
INV_X1 i_1_247 (.ZN (n_271), .A (n_1_143));
AOI222_X1 i_1_246 (.ZN (n_1_142), .A1 (n_1_169), .A2 (\m[5] ), .B1 (n_133), .B2 (hfn_ipo_n25)
    , .C1 (n_304), .C2 (hfn_ipo_n27));
INV_X1 i_1_245 (.ZN (n_270), .A (n_1_142));
AOI222_X1 i_1_244 (.ZN (n_1_141), .A1 (n_1_169), .A2 (\m[4] ), .B1 (n_132), .B2 (hfn_ipo_n25)
    , .C1 (n_303), .C2 (hfn_ipo_n27));
INV_X1 i_1_243 (.ZN (n_269), .A (n_1_141));
AOI222_X1 i_1_242 (.ZN (n_1_140), .A1 (n_1_169), .A2 (\m[3] ), .B1 (n_131), .B2 (hfn_ipo_n25)
    , .C1 (n_302), .C2 (hfn_ipo_n27));
INV_X1 i_1_241 (.ZN (n_268), .A (n_1_140));
AOI222_X1 i_1_240 (.ZN (n_1_139), .A1 (n_1_169), .A2 (\m[2] ), .B1 (n_130), .B2 (hfn_ipo_n25)
    , .C1 (n_301), .C2 (hfn_ipo_n27));
INV_X1 i_1_239 (.ZN (n_267), .A (n_1_139));
AOI222_X1 i_1_238 (.ZN (n_1_138), .A1 (n_1_169), .A2 (\m[1] ), .B1 (n_129), .B2 (hfn_ipo_n25)
    , .C1 (n_300), .C2 (hfn_ipo_n27));
INV_X1 i_1_237 (.ZN (n_266), .A (n_1_138));
AOI222_X1 i_1_236 (.ZN (n_1_137), .A1 (n_128), .A2 (hfn_ipo_n25), .B1 (n_1_169), .B2 (in1[0])
    , .C1 (hfn_ipo_n27), .C2 (n_299));
INV_X1 i_1_235 (.ZN (n_265), .A (n_1_137));
MUX2_X1 i_1_234 (.Z (n_1_136), .A (\res[31] ), .B (n_127), .S (n_1_174));
AND2_X2 i_1_229 (.ZN (n_1_135), .A1 (in2[31]), .A2 (n_1_170));
AOI22_X1 i_1_232 (.ZN (n_1_134), .A1 (n_1_180), .A2 (n_1_136), .B1 (n_1_135), .B2 (n_33));
INV_X1 i_1_231 (.ZN (n_264), .A (n_1_134));
AOI22_X1 i_1_230 (.ZN (n_1_133), .A1 (\res[30] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_126));
NOR4_X1 i_1_157 (.ZN (n_1_132), .A1 (n_1_182), .A2 (in2[31]), .A3 (resetReg), .A4 (reset));
AOI22_X1 i_1_228 (.ZN (n_1_131), .A1 (n_32), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[30]));
NAND2_X1 i_1_227 (.ZN (n_263), .A1 (n_1_131), .A2 (n_1_133));
AOI22_X1 i_1_226 (.ZN (n_1_130), .A1 (\res[29] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_125));
AOI22_X1 i_1_225 (.ZN (n_1_129), .A1 (n_31), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[29]));
NAND2_X1 i_1_224 (.ZN (n_262), .A1 (n_1_129), .A2 (n_1_130));
AOI22_X1 i_1_223 (.ZN (n_1_128), .A1 (\res[28] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_124));
AOI22_X1 i_1_222 (.ZN (n_1_127), .A1 (n_30), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[28]));
NAND2_X1 i_1_221 (.ZN (n_261), .A1 (n_1_127), .A2 (n_1_128));
AOI22_X1 i_1_220 (.ZN (n_1_126), .A1 (\res[27] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_123));
AOI22_X1 i_1_219 (.ZN (n_1_125), .A1 (n_29), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[27]));
NAND2_X1 i_1_218 (.ZN (n_260), .A1 (n_1_125), .A2 (n_1_126));
AOI22_X1 i_1_217 (.ZN (n_1_124), .A1 (\res[26] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_122));
AOI22_X1 i_1_216 (.ZN (n_1_123), .A1 (n_28), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[26]));
NAND2_X1 i_1_215 (.ZN (n_259), .A1 (n_1_123), .A2 (n_1_124));
AOI22_X1 i_1_214 (.ZN (n_1_122), .A1 (\res[25] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_121));
AOI22_X1 i_1_213 (.ZN (n_1_121), .A1 (n_27), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[25]));
NAND2_X1 i_1_212 (.ZN (n_258), .A1 (n_1_121), .A2 (n_1_122));
AOI22_X1 i_1_211 (.ZN (n_1_120), .A1 (\res[24] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_120));
AOI22_X1 i_1_210 (.ZN (n_1_119), .A1 (n_26), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[24]));
NAND2_X1 i_1_209 (.ZN (n_257), .A1 (n_1_119), .A2 (n_1_120));
AOI22_X1 i_1_208 (.ZN (n_1_118), .A1 (\res[23] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_119));
AOI22_X1 i_1_207 (.ZN (n_1_117), .A1 (n_25), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[23]));
NAND2_X1 i_1_206 (.ZN (n_256), .A1 (n_1_117), .A2 (n_1_118));
AOI22_X1 i_1_205 (.ZN (n_1_116), .A1 (\res[22] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_118));
AOI22_X1 i_1_204 (.ZN (n_1_115), .A1 (n_24), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[22]));
NAND2_X1 i_1_203 (.ZN (n_255), .A1 (n_1_115), .A2 (n_1_116));
AOI22_X1 i_1_202 (.ZN (n_1_114), .A1 (\res[21] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_117));
AOI22_X1 i_1_201 (.ZN (n_1_113), .A1 (n_23), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[21]));
NAND2_X1 i_1_200 (.ZN (n_254), .A1 (n_1_113), .A2 (n_1_114));
AOI22_X1 i_1_199 (.ZN (n_1_112), .A1 (\res[20] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_116));
AOI22_X1 i_1_198 (.ZN (n_1_111), .A1 (n_22), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[20]));
NAND2_X1 i_1_197 (.ZN (n_253), .A1 (n_1_111), .A2 (n_1_112));
AOI22_X1 i_1_196 (.ZN (n_1_110), .A1 (\res[19] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_115));
AOI22_X1 i_1_195 (.ZN (n_1_109), .A1 (n_21), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[19]));
NAND2_X1 i_1_194 (.ZN (n_252), .A1 (n_1_109), .A2 (n_1_110));
AOI22_X1 i_1_193 (.ZN (n_1_108), .A1 (\res[18] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_114));
AOI22_X1 i_1_192 (.ZN (n_1_107), .A1 (n_20), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[18]));
NAND2_X1 i_1_191 (.ZN (n_251), .A1 (n_1_107), .A2 (n_1_108));
AOI22_X1 i_1_190 (.ZN (n_1_106), .A1 (\res[17] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_113));
AOI22_X1 i_1_189 (.ZN (n_1_105), .A1 (n_19), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[17]));
NAND2_X1 i_1_188 (.ZN (n_250), .A1 (n_1_105), .A2 (n_1_106));
AOI22_X1 i_1_187 (.ZN (n_1_104), .A1 (\res[16] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_112));
AOI22_X1 i_1_186 (.ZN (n_1_103), .A1 (n_18), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[16]));
NAND2_X1 i_1_185 (.ZN (n_249), .A1 (n_1_103), .A2 (n_1_104));
AOI22_X1 i_1_184 (.ZN (n_1_102), .A1 (\res[15] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_111));
AOI22_X1 i_1_183 (.ZN (n_1_101), .A1 (n_17), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[15]));
NAND2_X1 i_1_182 (.ZN (n_248), .A1 (n_1_101), .A2 (n_1_102));
AOI22_X1 i_1_181 (.ZN (n_1_100), .A1 (\res[14] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_110));
AOI22_X1 i_1_180 (.ZN (n_1_99), .A1 (n_16), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[14]));
NAND2_X1 i_1_179 (.ZN (n_247), .A1 (n_1_99), .A2 (n_1_100));
AOI22_X1 i_1_178 (.ZN (n_1_98), .A1 (\res[13] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_109));
AOI22_X1 i_1_177 (.ZN (n_1_97), .A1 (n_15), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[13]));
NAND2_X1 i_1_176 (.ZN (n_246), .A1 (n_1_97), .A2 (n_1_98));
AOI22_X1 i_1_175 (.ZN (n_1_96), .A1 (\res[12] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_108));
AOI22_X1 i_1_174 (.ZN (n_1_95), .A1 (n_14), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[12]));
NAND2_X1 i_1_173 (.ZN (n_245), .A1 (n_1_95), .A2 (n_1_96));
AOI22_X1 i_1_172 (.ZN (n_1_94), .A1 (\res[11] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_107));
AOI22_X1 i_1_171 (.ZN (n_1_93), .A1 (n_13), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[11]));
NAND2_X1 i_1_170 (.ZN (n_244), .A1 (n_1_93), .A2 (n_1_94));
AOI22_X1 i_1_169 (.ZN (n_1_92), .A1 (\res[10] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_106));
AOI22_X1 i_1_168 (.ZN (n_1_91), .A1 (n_12), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[10]));
NAND2_X1 i_1_167 (.ZN (n_243), .A1 (n_1_91), .A2 (n_1_92));
AOI22_X1 i_1_166 (.ZN (n_1_90), .A1 (\res[9] ), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n25), .B2 (n_105));
AOI22_X1 i_1_165 (.ZN (n_1_89), .A1 (n_11), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[9]));
NAND2_X1 i_1_164 (.ZN (n_242), .A1 (n_1_89), .A2 (n_1_90));
AOI22_X1 i_1_163 (.ZN (n_1_88), .A1 (\res[8] ), .A2 (hfn_ipo_n28), .B1 (hfn_ipo_n26), .B2 (n_104));
AOI22_X1 i_1_162 (.ZN (n_1_87), .A1 (n_10), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[8]));
NAND2_X1 i_1_161 (.ZN (n_241), .A1 (n_1_87), .A2 (n_1_88));
AOI22_X1 i_1_160 (.ZN (n_1_86), .A1 (\res[7] ), .A2 (hfn_ipo_n28), .B1 (hfn_ipo_n26), .B2 (n_103));
AOI22_X1 i_1_159 (.ZN (n_1_85), .A1 (n_9), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[7]));
NAND2_X1 i_1_158 (.ZN (n_240), .A1 (n_1_85), .A2 (n_1_86));
AOI22_X1 i_1_156 (.ZN (n_1_84), .A1 (\res[6] ), .A2 (hfn_ipo_n28), .B1 (hfn_ipo_n26), .B2 (n_102));
AOI22_X1 i_1_155 (.ZN (n_1_83), .A1 (n_8), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[6]));
NAND2_X1 i_1_154 (.ZN (n_239), .A1 (n_1_83), .A2 (n_1_84));
AOI22_X1 i_1_153 (.ZN (n_1_81), .A1 (n_7), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[5]));
NAND2_X1 i_1_152 (.ZN (n_238), .A1 (n_1_81), .A2 (n_1_82));
AOI22_X1 i_1_151 (.ZN (n_1_80), .A1 (\res[4] ), .A2 (hfn_ipo_n28), .B1 (hfn_ipo_n26), .B2 (n_100));
AOI22_X1 i_1_150 (.ZN (n_1_79), .A1 (n_6), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[4]));
NAND2_X1 i_1_149 (.ZN (n_237), .A1 (n_1_79), .A2 (n_1_80));
AOI22_X1 i_1_148 (.ZN (n_1_78), .A1 (\res[3] ), .A2 (hfn_ipo_n28), .B1 (hfn_ipo_n26), .B2 (n_99));
AOI22_X1 i_1_147 (.ZN (n_1_77), .A1 (n_5), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[3]));
NAND2_X1 i_1_146 (.ZN (n_236), .A1 (n_1_77), .A2 (n_1_78));
AOI22_X1 i_1_145 (.ZN (n_1_76), .A1 (\res[2] ), .A2 (hfn_ipo_n28), .B1 (hfn_ipo_n26), .B2 (n_98));
AOI22_X1 i_1_144 (.ZN (n_1_75), .A1 (n_4), .A2 (n_1_135), .B1 (drc_ipo_n29), .B2 (in2[2]));
NAND2_X1 i_1_143 (.ZN (n_235), .A1 (n_1_75), .A2 (n_1_76));
AOI222_X1 i_1_142 (.ZN (n_1_74), .A1 (\res[1] ), .A2 (n_1_180), .B1 (n_1_135), .B2 (n_3)
    , .C1 (in2[1]), .C2 (drc_ipo_n29));
INV_X1 i_1_141 (.ZN (n_234), .A (n_1_74));
OAI22_X1 i_1_140 (.ZN (n_1_73), .A1 (en), .A2 (\counter[5] ), .B1 (n_335), .B2 (n_1_183));
AND2_X1 i_1_139 (.ZN (n_233), .A1 (n_1_178), .A2 (n_1_73));
AND2_X1 i_1_138 (.ZN (n_232), .A1 (n_1_73), .A2 (n_1_6));
AND2_X1 i_1_137 (.ZN (n_231), .A1 (n_1_73), .A2 (n_1_5));
AND2_X1 i_1_136 (.ZN (n_230), .A1 (n_1_73), .A2 (n_1_4));
AND2_X1 i_1_135 (.ZN (n_229), .A1 (n_1_73), .A2 (n_1_3));
AOI211_X1 i_1_134 (.ZN (n_228), .A (\counter[0] ), .B (n_335), .C1 (n_1_186), .C2 (\counter[5] ));
AND2_X1 i_1_133 (.ZN (n_1_72), .A1 (n_1_175), .A2 (n_1_184));
NOR2_X1 i_1_132 (.ZN (n_1_71), .A1 (n_335), .A2 (n_1_175));
AOI22_X1 i_1_131 (.ZN (n_1_70), .A1 (n_331), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_160));
INV_X1 i_1_130 (.ZN (n_227), .A (n_1_70));
AOI22_X1 i_1_129 (.ZN (n_1_69), .A1 (n_330), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_159));
INV_X1 i_1_128 (.ZN (n_226), .A (n_1_69));
AOI22_X1 i_1_127 (.ZN (n_1_68), .A1 (n_329), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_158));
INV_X1 i_1_126 (.ZN (n_225), .A (n_1_68));
AOI22_X1 i_1_125 (.ZN (n_1_67), .A1 (n_328), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_157));
INV_X1 i_1_124 (.ZN (n_224), .A (n_1_67));
AOI22_X1 i_1_123 (.ZN (n_1_66), .A1 (n_327), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_156));
INV_X1 i_1_122 (.ZN (n_223), .A (n_1_66));
AOI22_X1 i_1_121 (.ZN (n_1_65), .A1 (n_326), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_155));
INV_X1 i_1_120 (.ZN (n_222), .A (n_1_65));
AOI22_X1 i_1_119 (.ZN (n_1_64), .A1 (n_325), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_154));
INV_X1 i_1_118 (.ZN (n_221), .A (n_1_64));
AOI22_X1 i_1_117 (.ZN (n_1_63), .A1 (n_324), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_153));
INV_X1 i_1_116 (.ZN (n_220), .A (n_1_63));
AOI22_X1 i_1_115 (.ZN (n_1_62), .A1 (n_323), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_152));
INV_X1 i_1_114 (.ZN (n_219), .A (n_1_62));
AOI22_X1 i_1_113 (.ZN (n_1_61), .A1 (n_322), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_151));
INV_X1 i_1_112 (.ZN (n_218), .A (n_1_61));
AOI22_X1 i_1_111 (.ZN (n_1_60), .A1 (n_321), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_150));
INV_X1 i_1_110 (.ZN (n_217), .A (n_1_60));
AOI22_X1 i_1_109 (.ZN (n_1_59), .A1 (n_320), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_149));
INV_X1 i_1_108 (.ZN (n_216), .A (n_1_59));
AOI22_X1 i_1_107 (.ZN (n_1_58), .A1 (n_319), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_148));
INV_X1 i_1_106 (.ZN (n_215), .A (n_1_58));
AOI22_X1 i_1_105 (.ZN (n_1_57), .A1 (n_318), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_147));
INV_X1 i_1_104 (.ZN (n_214), .A (n_1_57));
AOI22_X1 i_1_103 (.ZN (n_1_56), .A1 (n_317), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_146));
INV_X1 i_1_102 (.ZN (n_213), .A (n_1_56));
AOI22_X1 i_1_101 (.ZN (n_1_55), .A1 (n_316), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_145));
INV_X1 i_1_100 (.ZN (n_212), .A (n_1_55));
AOI22_X1 i_1_99 (.ZN (n_1_54), .A1 (n_315), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_144));
INV_X1 i_1_98 (.ZN (n_211), .A (n_1_54));
AOI22_X1 i_1_97 (.ZN (n_1_53), .A1 (n_314), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_143));
INV_X1 i_1_96 (.ZN (n_210), .A (n_1_53));
AOI22_X1 i_1_95 (.ZN (n_1_52), .A1 (n_313), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_142));
INV_X1 i_1_94 (.ZN (n_209), .A (n_1_52));
AOI22_X1 i_1_93 (.ZN (n_1_51), .A1 (n_312), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_141));
INV_X1 i_1_92 (.ZN (n_208), .A (n_1_51));
AOI22_X1 i_1_91 (.ZN (n_1_50), .A1 (n_311), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_140));
INV_X1 i_1_90 (.ZN (n_207), .A (n_1_50));
AOI22_X1 i_1_89 (.ZN (n_1_49), .A1 (n_310), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_139));
INV_X1 i_1_88 (.ZN (n_206), .A (n_1_49));
AOI22_X1 i_1_87 (.ZN (n_1_48), .A1 (n_309), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_138));
INV_X1 i_1_86 (.ZN (n_205), .A (n_1_48));
AOI22_X1 i_1_85 (.ZN (n_1_47), .A1 (n_308), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_137));
INV_X1 i_1_84 (.ZN (n_204), .A (n_1_47));
AOI22_X1 i_1_83 (.ZN (n_1_46), .A1 (n_307), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_136));
INV_X1 i_1_82 (.ZN (n_203), .A (n_1_46));
AOI22_X1 i_1_81 (.ZN (n_1_45), .A1 (n_306), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_135));
INV_X1 i_1_80 (.ZN (n_202), .A (n_1_45));
AOI22_X1 i_1_79 (.ZN (n_1_44), .A1 (n_305), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_134));
INV_X1 i_1_78 (.ZN (n_201), .A (n_1_44));
AOI22_X1 i_1_77 (.ZN (n_1_43), .A1 (n_304), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_133));
INV_X1 i_1_76 (.ZN (n_200), .A (n_1_43));
AOI22_X1 i_1_75 (.ZN (n_1_42), .A1 (n_303), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_132));
INV_X1 i_1_74 (.ZN (n_199), .A (n_1_42));
AOI22_X1 i_1_73 (.ZN (n_1_41), .A1 (n_302), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_131));
INV_X1 i_1_72 (.ZN (n_198), .A (n_1_41));
AOI22_X1 i_1_71 (.ZN (n_1_40), .A1 (n_301), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_130));
INV_X1 i_1_70 (.ZN (n_197), .A (n_1_40));
AOI22_X1 i_1_69 (.ZN (n_1_39), .A1 (n_300), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_129));
INV_X1 i_1_68 (.ZN (n_196), .A (n_1_39));
AOI22_X1 i_1_67 (.ZN (n_1_38), .A1 (n_299), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_128));
INV_X1 i_1_66 (.ZN (n_195), .A (n_1_38));
AOI22_X1 i_1_65 (.ZN (n_1_37), .A1 (\res[31] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_127));
INV_X1 i_1_64 (.ZN (n_194), .A (n_1_37));
AOI22_X1 i_1_63 (.ZN (n_1_36), .A1 (\res[30] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_126));
INV_X1 i_1_62 (.ZN (n_193), .A (n_1_36));
AOI22_X1 i_1_61 (.ZN (n_1_35), .A1 (\res[29] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_125));
INV_X1 i_1_60 (.ZN (n_192), .A (n_1_35));
AOI22_X1 i_1_59 (.ZN (n_1_34), .A1 (\res[28] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_124));
INV_X1 i_1_58 (.ZN (n_191), .A (n_1_34));
AOI22_X1 i_1_57 (.ZN (n_1_33), .A1 (\res[27] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_123));
INV_X1 i_1_56 (.ZN (n_190), .A (n_1_33));
AOI22_X1 i_1_55 (.ZN (n_1_32), .A1 (\res[26] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_122));
INV_X1 i_1_54 (.ZN (n_189), .A (n_1_32));
AOI22_X1 i_1_53 (.ZN (n_1_31), .A1 (\res[25] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_121));
INV_X1 i_1_52 (.ZN (n_188), .A (n_1_31));
AOI22_X1 i_1_51 (.ZN (n_1_30), .A1 (\res[24] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_120));
INV_X1 i_1_50 (.ZN (n_187), .A (n_1_30));
AOI22_X1 i_1_49 (.ZN (n_1_29), .A1 (\res[23] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_119));
INV_X1 i_1_48 (.ZN (n_186), .A (n_1_29));
AOI22_X1 i_1_47 (.ZN (n_1_28), .A1 (\res[22] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_118));
INV_X1 i_1_46 (.ZN (n_185), .A (n_1_28));
AOI22_X1 i_1_45 (.ZN (n_1_27), .A1 (\res[21] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_117));
INV_X1 i_1_44 (.ZN (n_184), .A (n_1_27));
AOI22_X1 i_1_43 (.ZN (n_1_26), .A1 (\res[20] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_116));
INV_X1 i_1_42 (.ZN (n_183), .A (n_1_26));
AOI22_X1 i_1_41 (.ZN (n_1_25), .A1 (\res[19] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_115));
INV_X1 i_1_40 (.ZN (n_182), .A (n_1_25));
AOI22_X1 i_1_39 (.ZN (n_1_24), .A1 (\res[18] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_114));
INV_X1 i_1_38 (.ZN (n_181), .A (n_1_24));
AOI22_X1 i_1_37 (.ZN (n_1_23), .A1 (\res[17] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_113));
INV_X1 i_1_36 (.ZN (n_180), .A (n_1_23));
AOI22_X1 i_1_35 (.ZN (n_1_22), .A1 (\res[16] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_112));
INV_X1 i_1_34 (.ZN (n_179), .A (n_1_22));
AOI22_X1 i_1_33 (.ZN (n_1_21), .A1 (\res[15] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_111));
INV_X1 i_1_32 (.ZN (n_178), .A (n_1_21));
AOI22_X1 i_1_31 (.ZN (n_1_20), .A1 (\res[14] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_110));
INV_X1 i_1_30 (.ZN (n_177), .A (n_1_20));
AOI22_X1 i_1_29 (.ZN (n_1_19), .A1 (\res[13] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_109));
INV_X1 i_1_28 (.ZN (n_176), .A (n_1_19));
AOI22_X1 i_1_27 (.ZN (n_1_18), .A1 (\res[12] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_108));
INV_X1 i_1_26 (.ZN (n_175), .A (n_1_18));
AOI22_X1 i_1_25 (.ZN (n_1_17), .A1 (\res[11] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_107));
INV_X1 i_1_24 (.ZN (n_174), .A (n_1_17));
AOI22_X1 i_1_23 (.ZN (n_1_16), .A1 (\res[10] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_106));
INV_X1 i_1_22 (.ZN (n_173), .A (n_1_16));
AOI22_X1 i_1_21 (.ZN (n_1_15), .A1 (\res[9] ), .A2 (hfn_ipo_n23), .B1 (hfn_ipo_n21), .B2 (n_105));
INV_X1 i_1_20 (.ZN (n_172), .A (n_1_15));
AOI22_X1 i_1_19 (.ZN (n_1_14), .A1 (\res[8] ), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_104));
INV_X1 i_1_18 (.ZN (n_171), .A (n_1_14));
AOI22_X1 i_1_17 (.ZN (n_1_13), .A1 (\res[7] ), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_103));
INV_X1 i_1_16 (.ZN (n_170), .A (n_1_13));
AOI22_X1 i_1_15 (.ZN (n_1_12), .A1 (\res[6] ), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_102));
INV_X1 i_1_14 (.ZN (n_169), .A (n_1_12));
AOI22_X1 i_1_13 (.ZN (n_1_11), .A1 (\res[5] ), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_101));
INV_X1 i_1_12 (.ZN (n_168), .A (n_1_11));
AOI22_X1 i_1_11 (.ZN (n_1_10), .A1 (\res[4] ), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_100));
INV_X1 i_1_10 (.ZN (n_167), .A (n_1_10));
AOI22_X1 i_1_9 (.ZN (n_1_9), .A1 (\res[3] ), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_99));
INV_X1 i_1_8 (.ZN (n_166), .A (n_1_9));
AOI22_X1 i_1_7 (.ZN (n_1_8), .A1 (\res[2] ), .A2 (hfn_ipo_n24), .B1 (hfn_ipo_n22), .B2 (n_98));
INV_X1 i_1_6 (.ZN (n_165), .A (n_1_8));
AND2_X1 i_1_5 (.ZN (n_164), .A1 (n_1_184), .A2 (\res[1] ));
AND2_X1 i_1_4 (.ZN (n_163), .A1 (en), .A2 (reset));
HA_X1 i_1_3 (.CO (n_1_7), .S (n_1_6), .A (\counter[4] ), .B (n_1_2));
HA_X1 i_1_2 (.CO (n_1_2), .S (n_1_5), .A (\counter[3] ), .B (n_1_1));
HA_X1 i_1_1 (.CO (n_1_1), .S (n_1_4), .A (\counter[2] ), .B (n_1_0));
HA_X1 i_1_0 (.CO (n_1_0), .S (n_1_3), .A (\counter[1] ), .B (\counter[0] ));
DFF_X1 \res_reg[0]  (.Q (\res[0] ), .CK (CTS_n_tid1_32), .D (n_234));
DFF_X1 \res_reg[1]  (.Q (\res[1] ), .CK (CTS_n_tid1_33), .D (n_235));
DFF_X1 \res_reg[2]  (.Q (\res[2] ), .CK (CTS_n_tid1_33), .D (n_236));
DFF_X1 \res_reg[3]  (.Q (\res[3] ), .CK (CTS_n_tid1_33), .D (n_237));
DFF_X1 \res_reg[4]  (.Q (\res[4] ), .CK (CTS_n_tid1_33), .D (n_238));
DFF_X1 \res_reg[5]  (.Q (\res[5] ), .CK (CTS_n_tid1_33), .D (n_239));
DFF_X1 \res_reg[6]  (.Q (\res[6] ), .CK (CTS_n_tid1_33), .D (n_240));
DFF_X1 \res_reg[7]  (.Q (\res[7] ), .CK (CTS_n_tid1_33), .D (n_241));
DFF_X1 \res_reg[8]  (.Q (\res[8] ), .CK (CTS_n_tid1_33), .D (n_242));
DFF_X1 \res_reg[9]  (.Q (\res[9] ), .CK (CTS_n_tid1_32), .D (n_243));
DFF_X1 \res_reg[10]  (.Q (\res[10] ), .CK (CTS_n_tid1_32), .D (n_244));
DFF_X1 \res_reg[11]  (.Q (\res[11] ), .CK (CTS_n_tid1_32), .D (n_245));
DFF_X1 \res_reg[12]  (.Q (\res[12] ), .CK (CTS_n_tid1_32), .D (n_246));
DFF_X1 \res_reg[13]  (.Q (\res[13] ), .CK (CTS_n_tid1_32), .D (n_247));
DFF_X1 \res_reg[14]  (.Q (\res[14] ), .CK (CTS_n_tid1_32), .D (n_248));
DFF_X1 \res_reg[15]  (.Q (\res[15] ), .CK (CTS_n_tid1_32), .D (n_249));
DFF_X1 \res_reg[16]  (.Q (\res[16] ), .CK (CTS_n_tid1_32), .D (n_250));
DFF_X1 \res_reg[17]  (.Q (\res[17] ), .CK (CTS_n_tid1_32), .D (n_251));
DFF_X1 \res_reg[18]  (.Q (\res[18] ), .CK (CTS_n_tid1_32), .D (n_252));
DFF_X1 \res_reg[19]  (.Q (\res[19] ), .CK (CTS_n_tid1_32), .D (n_253));
DFF_X1 \res_reg[20]  (.Q (\res[20] ), .CK (CTS_n_tid1_32), .D (n_254));
DFF_X1 \res_reg[21]  (.Q (\res[21] ), .CK (CTS_n_tid1_32), .D (n_255));
DFF_X1 \res_reg[22]  (.Q (\res[22] ), .CK (CTS_n_tid1_32), .D (n_256));
DFF_X1 \res_reg[23]  (.Q (\res[23] ), .CK (CTS_n_tid1_32), .D (n_257));
DFF_X1 \res_reg[24]  (.Q (\res[24] ), .CK (CTS_n_tid1_32), .D (n_258));
DFF_X1 \res_reg[25]  (.Q (\res[25] ), .CK (CTS_n_tid1_32), .D (n_259));
DFF_X1 \res_reg[26]  (.Q (\res[26] ), .CK (CTS_n_tid1_32), .D (n_260));
DFF_X1 \res_reg[27]  (.Q (\res[27] ), .CK (CTS_n_tid1_32), .D (n_261));
DFF_X1 \res_reg[28]  (.Q (\res[28] ), .CK (CTS_n_tid1_32), .D (n_262));
DFF_X1 \res_reg[29]  (.Q (\res[29] ), .CK (CTS_n_tid1_32), .D (n_263));
DFF_X1 \res_reg[30]  (.Q (\res[30] ), .CK (CTS_n_tid1_32), .D (n_264));
DFF_X1 \res_reg[31]  (.Q (\res[31] ), .CK (CTS_n_tid1_32), .D (n_265));
DFF_X1 \res_reg[32]  (.Q (\res[32] ), .CK (CTS_n_tid1_32), .D (n_266));
DFF_X1 \res_reg[33]  (.Q (\res[33] ), .CK (CTS_n_tid1_32), .D (n_267));
DFF_X1 \res_reg[34]  (.Q (\res[34] ), .CK (CTS_n_tid1_32), .D (n_268));
DFF_X1 \res_reg[35]  (.Q (\res[35] ), .CK (CTS_n_tid1_32), .D (n_269));
DFF_X1 \res_reg[36]  (.Q (\res[36] ), .CK (CTS_n_tid1_32), .D (n_270));
DFF_X1 \res_reg[37]  (.Q (\res[37] ), .CK (CTS_n_tid1_32), .D (n_271));
DFF_X1 \res_reg[38]  (.Q (\res[38] ), .CK (CTS_n_tid1_32), .D (n_272));
DFF_X1 \res_reg[39]  (.Q (\res[39] ), .CK (CTS_n_tid1_32), .D (n_273));
DFF_X1 \res_reg[40]  (.Q (\res[40] ), .CK (CTS_n_tid1_32), .D (n_274));
DFF_X1 \res_reg[41]  (.Q (\res[41] ), .CK (CTS_n_tid1_33), .D (n_275));
DFF_X1 \res_reg[42]  (.Q (\res[42] ), .CK (CTS_n_tid1_33), .D (n_276));
DFF_X1 \res_reg[43]  (.Q (\res[43] ), .CK (CTS_n_tid1_33), .D (n_277));
DFF_X1 \res_reg[44]  (.Q (\res[44] ), .CK (CTS_n_tid1_33), .D (n_278));
DFF_X1 \res_reg[45]  (.Q (\res[45] ), .CK (CTS_n_tid1_33), .D (n_279));
DFF_X1 \res_reg[46]  (.Q (\res[46] ), .CK (CTS_n_tid1_33), .D (n_280));
DFF_X1 \res_reg[47]  (.Q (\res[47] ), .CK (CTS_n_tid1_33), .D (n_281));
DFF_X1 \res_reg[48]  (.Q (\res[48] ), .CK (CTS_n_tid1_33), .D (n_282));
DFF_X1 \res_reg[49]  (.Q (\res[49] ), .CK (CTS_n_tid1_33), .D (n_283));
DFF_X1 \res_reg[50]  (.Q (\res[50] ), .CK (CTS_n_tid1_33), .D (n_284));
DFF_X1 \res_reg[51]  (.Q (\res[51] ), .CK (CTS_n_tid1_33), .D (n_285));
DFF_X1 \res_reg[52]  (.Q (\res[52] ), .CK (CTS_n_tid1_33), .D (n_286));
DFF_X1 \res_reg[53]  (.Q (\res[53] ), .CK (CTS_n_tid1_33), .D (n_287));
DFF_X1 \res_reg[54]  (.Q (\res[54] ), .CK (CTS_n_tid1_33), .D (n_288));
DFF_X1 \res_reg[55]  (.Q (\res[55] ), .CK (CTS_n_tid1_33), .D (n_289));
DFF_X1 \res_reg[56]  (.Q (\res[56] ), .CK (CTS_n_tid1_33), .D (n_290));
DFF_X1 \res_reg[57]  (.Q (\res[57] ), .CK (CTS_n_tid1_33), .D (n_291));
DFF_X1 \res_reg[58]  (.Q (\res[58] ), .CK (CTS_n_tid1_33), .D (n_292));
DFF_X1 \res_reg[59]  (.Q (\res[59] ), .CK (CTS_n_tid1_33), .D (n_293));
DFF_X1 \res_reg[60]  (.Q (\res[60] ), .CK (CTS_n_tid1_33), .D (n_294));
DFF_X1 \res_reg[61]  (.Q (\res[61] ), .CK (CTS_n_tid1_33), .D (n_295));
DFF_X1 \res_reg[62]  (.Q (\res[62] ), .CK (CTS_n_tid1_33), .D (n_296));
DFF_X1 \res_reg[63]  (.Q (\res[63] ), .CK (CTS_n_tid1_33), .D (n_297));
DFF_X1 \res_reg[64]  (.Q (\res[64] ), .CK (CTS_n_tid1_33), .D (n_298));
CLKGATETST_X8 clk_gate_res_reg (.GCK (CTS_n_tid1_82), .CK (clk_CTS_0_PP_1), .E (n_332), .SE (1'b0 ));
MUX2_X1 resetReg_reg_enable_mux_0 (.Z (n_162), .A (resetReg), .B (n_163), .S (n_335));
DFF_X1 resetReg_reg (.Q (resetReg), .CK (CTS_n_tid0_179), .D (n_162));
DFF_X1 \counter_reg[0]  (.Q (\counter[0] ), .CK (n_1), .D (n_228));
DFF_X1 \counter_reg[1]  (.Q (\counter[1] ), .CK (n_1), .D (n_229));
DFF_X1 \counter_reg[2]  (.Q (\counter[2] ), .CK (n_1), .D (n_230));
DFF_X1 \counter_reg[3]  (.Q (\counter[3] ), .CK (n_1), .D (n_231));
DFF_X1 \counter_reg[4]  (.Q (\counter[4] ), .CK (n_1), .D (n_232));
DFF_X1 \counter_reg[5]  (.Q (\counter[5] ), .CK (n_1), .D (n_233));
CLKGATETST_X1 clk_gate_counter_reg (.GCK (n_1), .CK (clk_CTS_0_PP_0), .E (en), .SE (1'b0 ));
DFF_X1 \result_reg[0]  (.Q (result[0]), .CK (CTS_n_tid0_91), .D (n_164));
DFF_X1 \result_reg[1]  (.Q (result[1]), .CK (CTS_n_tid0_91), .D (n_165));
DFF_X1 \result_reg[2]  (.Q (result[2]), .CK (CTS_n_tid0_91), .D (n_166));
DFF_X1 \result_reg[3]  (.Q (result[3]), .CK (CTS_n_tid0_91), .D (n_167));
DFF_X1 \result_reg[4]  (.Q (result[4]), .CK (CTS_n_tid0_91), .D (n_168));
DFF_X1 \result_reg[5]  (.Q (result[5]), .CK (CTS_n_tid0_91), .D (n_169));
DFF_X1 \result_reg[6]  (.Q (result[6]), .CK (CTS_n_tid0_91), .D (n_170));
DFF_X1 \result_reg[7]  (.Q (result[7]), .CK (CTS_n_tid0_91), .D (n_171));
DFF_X1 \result_reg[8]  (.Q (result[8]), .CK (CTS_n_tid0_91), .D (n_172));
DFF_X1 \result_reg[9]  (.Q (result[9]), .CK (CTS_n_tid0_91), .D (n_173));
DFF_X1 \result_reg[10]  (.Q (result[10]), .CK (CTS_n_tid0_91), .D (n_174));
DFF_X1 \result_reg[11]  (.Q (result[11]), .CK (CTS_n_tid0_91), .D (n_175));
DFF_X1 \result_reg[12]  (.Q (result[12]), .CK (CTS_n_tid0_91), .D (n_176));
DFF_X1 \result_reg[13]  (.Q (result[13]), .CK (CTS_n_tid0_91), .D (n_177));
DFF_X1 \result_reg[14]  (.Q (result[14]), .CK (CTS_n_tid0_91), .D (n_178));
DFF_X1 \result_reg[15]  (.Q (result[15]), .CK (CTS_n_tid0_91), .D (n_179));
DFF_X1 \result_reg[16]  (.Q (result[16]), .CK (CTS_n_tid0_91), .D (n_180));
DFF_X1 \result_reg[17]  (.Q (result[17]), .CK (CTS_n_tid0_91), .D (n_181));
DFF_X1 \result_reg[18]  (.Q (result[18]), .CK (CTS_n_tid0_91), .D (n_182));
DFF_X1 \result_reg[19]  (.Q (result[19]), .CK (CTS_n_tid0_91), .D (n_183));
DFF_X1 \result_reg[20]  (.Q (result[20]), .CK (CTS_n_tid0_91), .D (n_184));
DFF_X1 \result_reg[21]  (.Q (result[21]), .CK (CTS_n_tid0_91), .D (n_185));
DFF_X1 \result_reg[22]  (.Q (result[22]), .CK (CTS_n_tid0_91), .D (n_186));
DFF_X1 \result_reg[23]  (.Q (result[23]), .CK (CTS_n_tid0_91), .D (n_187));
DFF_X1 \result_reg[24]  (.Q (result[24]), .CK (CTS_n_tid0_91), .D (n_188));
DFF_X1 \result_reg[25]  (.Q (result[25]), .CK (CTS_n_tid0_91), .D (n_189));
DFF_X1 \result_reg[26]  (.Q (result[26]), .CK (CTS_n_tid0_91), .D (n_190));
DFF_X1 \result_reg[27]  (.Q (result[27]), .CK (CTS_n_tid0_91), .D (n_191));
DFF_X1 \result_reg[28]  (.Q (result[28]), .CK (CTS_n_tid0_91), .D (n_192));
DFF_X1 \result_reg[29]  (.Q (result[29]), .CK (CTS_n_tid0_91), .D (n_193));
DFF_X1 \result_reg[30]  (.Q (result[30]), .CK (CTS_n_tid0_91), .D (n_194));
DFF_X1 \result_reg[31]  (.Q (result[31]), .CK (CTS_n_tid0_91), .D (n_195));
DFF_X1 \result_reg[32]  (.Q (result[32]), .CK (CTS_n_tid0_91), .D (n_196));
DFF_X1 \result_reg[33]  (.Q (result[33]), .CK (CTS_n_tid0_91), .D (n_197));
DFF_X1 \result_reg[34]  (.Q (result[34]), .CK (CTS_n_tid0_91), .D (n_198));
DFF_X1 \result_reg[35]  (.Q (result[35]), .CK (CTS_n_tid0_91), .D (n_199));
DFF_X1 \result_reg[36]  (.Q (result[36]), .CK (CTS_n_tid0_91), .D (n_200));
DFF_X1 \result_reg[37]  (.Q (result[37]), .CK (CTS_n_tid0_91), .D (n_201));
DFF_X1 \result_reg[38]  (.Q (result[38]), .CK (CTS_n_tid0_91), .D (n_202));
DFF_X1 \result_reg[39]  (.Q (result[39]), .CK (CTS_n_tid0_91), .D (n_203));
DFF_X1 \result_reg[40]  (.Q (result[40]), .CK (CTS_n_tid0_91), .D (n_204));
DFF_X1 \result_reg[41]  (.Q (result[41]), .CK (CTS_n_tid0_91), .D (n_205));
DFF_X1 \result_reg[42]  (.Q (result[42]), .CK (CTS_n_tid0_91), .D (n_206));
DFF_X1 \result_reg[43]  (.Q (result[43]), .CK (CTS_n_tid0_91), .D (n_207));
DFF_X1 \result_reg[44]  (.Q (result[44]), .CK (CTS_n_tid0_91), .D (n_208));
DFF_X1 \result_reg[45]  (.Q (result[45]), .CK (CTS_n_tid0_91), .D (n_209));
DFF_X1 \result_reg[46]  (.Q (result[46]), .CK (CTS_n_tid0_91), .D (n_210));
DFF_X1 \result_reg[47]  (.Q (result[47]), .CK (CTS_n_tid0_91), .D (n_211));
DFF_X1 \result_reg[48]  (.Q (result[48]), .CK (CTS_n_tid0_91), .D (n_212));
DFF_X1 \result_reg[49]  (.Q (result[49]), .CK (CTS_n_tid0_91), .D (n_213));
DFF_X1 \result_reg[50]  (.Q (result[50]), .CK (CTS_n_tid0_91), .D (n_214));
DFF_X1 \result_reg[51]  (.Q (result[51]), .CK (CTS_n_tid0_91), .D (n_215));
DFF_X1 \result_reg[52]  (.Q (result[52]), .CK (CTS_n_tid0_91), .D (n_216));
DFF_X1 \result_reg[53]  (.Q (result[53]), .CK (CTS_n_tid0_91), .D (n_217));
DFF_X1 \result_reg[54]  (.Q (result[54]), .CK (CTS_n_tid0_91), .D (n_218));
DFF_X1 \result_reg[55]  (.Q (result[55]), .CK (CTS_n_tid0_91), .D (n_219));
DFF_X1 \result_reg[56]  (.Q (result[56]), .CK (CTS_n_tid0_91), .D (n_220));
DFF_X1 \result_reg[57]  (.Q (result[57]), .CK (CTS_n_tid0_91), .D (n_221));
DFF_X1 \result_reg[58]  (.Q (result[58]), .CK (CTS_n_tid0_91), .D (n_222));
DFF_X1 \result_reg[59]  (.Q (result[59]), .CK (CTS_n_tid0_91), .D (n_223));
DFF_X1 \result_reg[60]  (.Q (result[60]), .CK (CTS_n_tid0_91), .D (n_224));
DFF_X1 \result_reg[61]  (.Q (result[61]), .CK (CTS_n_tid0_91), .D (n_225));
DFF_X1 \result_reg[62]  (.Q (result[62]), .CK (CTS_n_tid0_91), .D (n_226));
DFF_X1 \result_reg[63]  (.Q (result[63]), .CK (CTS_n_tid0_91), .D (n_227));
CLKGATETST_X4 clk_gate_result_reg (.GCK (CTS_n_tid0_92), .CK (clk_CTS_0_PP_15), .E (n_333), .SE (1'b0 ));
datapath__0_11 i_11 (.p_0 ({n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, 
    n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, 
    n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, 
    n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, n_121, 
    n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, 
    n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
    uc_2}), .p_1 ({1'b0 , n_331, n_330, n_329, n_328, n_327, n_326, n_325, n_324, 
    n_323, n_322, n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314, n_313, 
    n_312, n_311, n_310, n_309, n_308, n_307, n_306, n_305, n_304, n_303, n_302, 
    n_301, n_300, n_299, \res[31] , \res[30] , \res[29] , \res[28] , \res[27] , \res[26] , 
    \res[25] , \res[24] , \res[23] , \res[22] , \res[21] , \res[20] , \res[19] , 
    \res[18] , \res[17] , \res[16] , \res[15] , \res[14] , \res[13] , \res[12] , 
    \res[11] , \res[10] , \res[9] , \res[8] , \res[7] , \res[6] , \res[5] , \res[4] , 
    \res[3] , \res[2] , \res[1] }));
datapath__0_9 i_9 (.p_1 ({n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, 
    n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, 
    n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65}), .m ({\m[31] , \m[30] , 
    \m[29] , \m[28] , \m[27] , \m[26] , \m[25] , \m[24] , \m[23] , \m[22] , \m[21] , 
    \m[20] , \m[19] , \m[18] , \m[17] , \m[16] , \m[15] , \m[14] , \m[13] , \m[12] , 
    \m[11] , \m[10] , \m[9] , \m[8] , \m[7] , \m[6] , \m[5] , \m[4] , \m[3] , \m[2] , 
    \m[1] , in1[0]}), .p_0 ({\res[63] , \res[62] , \res[61] , \res[60] , \res[59] , 
    \res[58] , \res[57] , \res[56] , \res[55] , \res[54] , \res[53] , \res[52] , 
    \res[51] , \res[50] , \res[49] , \res[48] , \res[47] , \res[46] , \res[45] , 
    \res[44] , \res[43] , \res[42] , \res[41] , \res[40] , \res[39] , \res[38] , 
    \res[37] , \res[36] , \res[35] , \res[34] , \res[33] , \res[32] }));
DFF_X1 enableOutput_reg (.Q (enableOutput), .CK (CTS_n_tid0_179), .D (n_334));
datapath__0_2 i_2 (.p_0 ({n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
    n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, uc_1}), .in1 ({in1[31], in1[30], 
    in1[29], in1[28], in1[27], in1[26], in1[25], in1[24], in1[23], in1[22], in1[21], 
    in1[20], in1[19], in1[18], in1[17], in1[16], in1[15], in1[14], in1[13], in1[12], 
    in1[11], in1[10], in1[9], in1[8], in1[7], in1[6], in1[5], in1[4], in1[3], in1[2], 
    in1[1], in1[0]}));
datapath i_0 (.p_0 ({n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
    n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, 
    n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, uc_0}), .in2 ({in2[31], in2[30], in2[29], 
    in2[28], in2[27], in2[26], in2[25], in2[24], in2[23], in2[22], in2[21], in2[20], 
    in2[19], in2[18], in2[17], in2[16], in2[15], in2[14], in2[13], in2[12], in2[11], 
    in2[10], in2[9], in2[8], in2[7], in2[6], in2[5], in2[4], in2[3], in2[2], in2[1], 
    in2[0]}));
CLKBUF_X2 hfn_ipo_c22 (.Z (hfn_ipo_n22), .A (n_1_71));
CLKBUF_X2 hfn_ipo_c23 (.Z (hfn_ipo_n23), .A (n_1_72));
CLKBUF_X2 hfn_ipo_c24 (.Z (hfn_ipo_n24), .A (n_1_72));
CLKBUF_X2 hfn_ipo_c25 (.Z (hfn_ipo_n25), .A (n_1_172));
CLKBUF_X2 hfn_ipo_c27 (.Z (hfn_ipo_n27), .A (n_1_173));
CLKBUF_X2 hfn_ipo_c28 (.Z (hfn_ipo_n28), .A (n_1_173));
CLKBUF_X2 drc_ipo_c29 (.Z (drc_ipo_n29), .A (n_1_132));
BUF_X4 drc_ipo_c30 (.Z (drc_ipo_n30), .A (\res[0] ));
CLKBUF_X2 hfn_ipo_c26 (.Z (hfn_ipo_n26), .A (n_1_172));
CLKBUF_X2 hfn_ipo_c21 (.Z (hfn_ipo_n21), .A (n_1_71));
CLKBUF_X3 CTS_L3_c_tid1_35 (.Z (CTS_n_tid1_32), .A (CTS_n_tid1_82));
CLKBUF_X3 CTS_L3_c_tid1_36 (.Z (CTS_n_tid1_33), .A (CTS_n_tid1_82));
CLKBUF_X3 CTS_L3_c_tid0_79 (.Z (CTS_n_tid0_91), .A (CTS_n_tid0_92));
CLKBUF_X1 CTS_L3_c_tid0_148 (.Z (CTS_n_tid0_179), .A (clk_CTS_0_PP_0));
CLKBUF_X1 CTS_L1_c_tid0_153 (.Z (clk_CTS_0_PP_1), .A (CTSclk_CTS_0_PP_15PP_0));

endmodule //sequentialmultiplier

module registerNbits__0_25 (clk_CTS_0_PP_11, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_11;
wire CLOCK_slh__n79;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CLOCK_slh__n83;
wire CLOCK_slh__n81;
wire CLOCK_slh__n85;
wire CLOCK_slh__n87;
wire CLOCK_slh__n89;
wire CLOCK_slh__n91;
wire CLOCK_slh__n93;
wire CLOCK_slh__n95;
wire CLOCK_slh__n97;
wire CLOCK_slh__n99;
wire CLOCK_slh__n101;
wire CLOCK_slh__n103;
wire CLOCK_slh__n105;
wire CLOCK_slh__n107;
wire CLOCK_slh__n109;
wire CLOCK_slh__n111;
wire CLOCK_slh__n113;
wire CLOCK_slh__n115;
wire CLOCK_slh__n117;
wire CLOCK_slh__n119;
wire CLOCK_slh__n121;
wire CLOCK_slh__n123;
wire CLOCK_slh__n125;
wire CLOCK_slh__n127;
wire CLOCK_slh__n129;
wire CLOCK_slh__n131;
wire CLOCK_slh__n133;
wire CLOCK_slh__n135;
wire CLOCK_slh__n137;
wire CLOCK_slh__n139;
wire CLOCK_slh__n141;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n141), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n137), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n135), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n111), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n99), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n129), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n97), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n131), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n113), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n121), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n109), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n95), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n93), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n91), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n89), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n115), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n87), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n85), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n123), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n127), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n133), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n83), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n81), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n79), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n119), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n117), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n103), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n101), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n125), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n107), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n105), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n139), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTS_0_PP_11), .E (n_1), .SE (1'b0 ));
CLKBUF_X1 CLOCK_slh__c41 (.Z (n_10), .A (CLOCK_slh__n79));
CLKBUF_X1 CLOCK_slh__c45 (.Z (n_12), .A (CLOCK_slh__n83));
CLKBUF_X1 CLOCK_slh__c43 (.Z (n_11), .A (CLOCK_slh__n81));
CLKBUF_X1 CLOCK_slh__c47 (.Z (n_16), .A (CLOCK_slh__n85));
CLKBUF_X1 CLOCK_slh__c49 (.Z (n_17), .A (CLOCK_slh__n87));
CLKBUF_X1 CLOCK_slh__c51 (.Z (n_19), .A (CLOCK_slh__n89));
CLKBUF_X1 CLOCK_slh__c53 (.Z (n_20), .A (CLOCK_slh__n91));
CLKBUF_X1 CLOCK_slh__c55 (.Z (n_21), .A (CLOCK_slh__n93));
CLKBUF_X1 CLOCK_slh__c57 (.Z (n_22), .A (CLOCK_slh__n95));
CLKBUF_X1 CLOCK_slh__c59 (.Z (n_27), .A (CLOCK_slh__n97));
CLKBUF_X1 CLOCK_slh__c61 (.Z (n_29), .A (CLOCK_slh__n99));
CLKBUF_X1 CLOCK_slh__c63 (.Z (n_6), .A (CLOCK_slh__n101));
CLKBUF_X1 CLOCK_slh__c65 (.Z (n_7), .A (CLOCK_slh__n103));
CLKBUF_X1 CLOCK_slh__c67 (.Z (n_3), .A (CLOCK_slh__n105));
CLKBUF_X1 CLOCK_slh__c69 (.Z (n_4), .A (CLOCK_slh__n107));
CLKBUF_X1 CLOCK_slh__c71 (.Z (n_23), .A (CLOCK_slh__n109));
CLKBUF_X1 CLOCK_slh__c73 (.Z (n_30), .A (CLOCK_slh__n111));
CLKBUF_X1 CLOCK_slh__c75 (.Z (n_25), .A (CLOCK_slh__n113));
CLKBUF_X1 CLOCK_slh__c77 (.Z (n_18), .A (CLOCK_slh__n115));
CLKBUF_X1 CLOCK_slh__c79 (.Z (n_8), .A (CLOCK_slh__n117));
CLKBUF_X1 CLOCK_slh__c81 (.Z (n_9), .A (CLOCK_slh__n119));
CLKBUF_X1 CLOCK_slh__c83 (.Z (n_24), .A (CLOCK_slh__n121));
CLKBUF_X1 CLOCK_slh__c85 (.Z (n_15), .A (CLOCK_slh__n123));
CLKBUF_X1 CLOCK_slh__c87 (.Z (n_5), .A (CLOCK_slh__n125));
CLKBUF_X1 CLOCK_slh__c89 (.Z (n_14), .A (CLOCK_slh__n127));
CLKBUF_X1 CLOCK_slh__c91 (.Z (n_28), .A (CLOCK_slh__n129));
CLKBUF_X1 CLOCK_slh__c93 (.Z (n_26), .A (CLOCK_slh__n131));
CLKBUF_X1 CLOCK_slh__c95 (.Z (n_13), .A (CLOCK_slh__n133));
CLKBUF_X1 CLOCK_slh__c97 (.Z (n_31), .A (CLOCK_slh__n135));
CLKBUF_X1 CLOCK_slh__c99 (.Z (n_32), .A (CLOCK_slh__n137));
CLKBUF_X1 CLOCK_slh__c101 (.Z (n_2), .A (CLOCK_slh__n139));
CLKBUF_X1 CLOCK_slh__c103 (.Z (n_33), .A (CLOCK_slh__n141));

endmodule //registerNbits__0_25

module registerNbits__0_22 (clk_CTS_0_PP_0, clk_CTS_0_PP_3, clk, reset, en, inp, 
    out);

output [31:0] out;
output clk_CTS_0_PP_0;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_3;
wire drc_ipo_n6;
wire n_0_0;
wire n_1;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid0_12;
wire CTS_n_tid0_13;
wire CTS_n_tid0_14;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid0_14), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid0_14), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid0_14), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid0_14), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid0_14), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid0_14), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid0_14), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid0_14), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid0_14), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid0_14), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid0_14), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid0_14), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid0_14), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid0_14), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid0_14), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid0_14), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid0_13), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid0_13), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid0_13), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid0_13), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid0_13), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid0_13), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid0_13), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid0_13), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid0_13), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid0_13), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid0_13), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid0_13), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid0_13), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid0_13), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid0_13), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n6), .CK (CTS_n_tid0_14), .D (n_33));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n_tid0_12), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
BUF_X4 drc_ipo_c3 (.Z (out[31]), .A (drc_ipo_n6));
CLKBUF_X1 CTS_L2_c_tid0_18 (.Z (clk_CTS_0_PP_0), .A (clk_CTS_0_PP_3));
CLKBUF_X3 CTS_L4_c_tid0_8 (.Z (CTS_n_tid0_13), .A (CTS_n_tid0_12));
CLKBUF_X3 CTS_L4_c_tid0_9 (.Z (CTS_n_tid0_14), .A (CTS_n_tid0_12));

endmodule //registerNbits__0_22

module integrationMult (inputA, inputB, clk, reset, en, result);

output [63:0] result;
input clk;
input en;
input [31:0] inputA;
input [31:0] inputB;
input reset;
wire CTS_n_tid0_3;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire enableOutput;
wire \outB_reg[31] ;
wire \outB_reg[30] ;
wire \outB_reg[29] ;
wire \outB_reg[28] ;
wire \outB_reg[27] ;
wire \outB_reg[26] ;
wire \outB_reg[25] ;
wire \outB_reg[24] ;
wire \outB_reg[23] ;
wire \outB_reg[22] ;
wire \outB_reg[21] ;
wire \outB_reg[20] ;
wire \outB_reg[19] ;
wire \outB_reg[18] ;
wire \outB_reg[17] ;
wire \outB_reg[16] ;
wire \outB_reg[15] ;
wire \outB_reg[14] ;
wire \outB_reg[13] ;
wire \outB_reg[12] ;
wire \outB_reg[11] ;
wire \outB_reg[10] ;
wire \outB_reg[9] ;
wire \outB_reg[8] ;
wire \outB_reg[7] ;
wire \outB_reg[6] ;
wire \outB_reg[5] ;
wire \outB_reg[4] ;
wire \outB_reg[3] ;
wire \outB_reg[2] ;
wire \outB_reg[1] ;
wire \outB_reg[0] ;
wire \outA_reg[31] ;
wire \outA_reg[30] ;
wire \outA_reg[29] ;
wire \outA_reg[28] ;
wire \outA_reg[27] ;
wire \outA_reg[26] ;
wire \outA_reg[25] ;
wire \outA_reg[24] ;
wire \outA_reg[23] ;
wire \outA_reg[22] ;
wire \outA_reg[21] ;
wire \outA_reg[20] ;
wire \outA_reg[19] ;
wire \outA_reg[18] ;
wire \outA_reg[17] ;
wire \outA_reg[16] ;
wire \outA_reg[15] ;
wire \outA_reg[14] ;
wire \outA_reg[13] ;
wire \outA_reg[12] ;
wire \outA_reg[11] ;
wire \outA_reg[10] ;
wire \outA_reg[9] ;
wire \outA_reg[8] ;
wire \outA_reg[7] ;
wire \outA_reg[6] ;
wire \outA_reg[5] ;
wire \outA_reg[4] ;
wire \outA_reg[3] ;
wire \outA_reg[2] ;
wire \outA_reg[1] ;
wire \outA_reg[0] ;
wire CTS_n_tid0_6;
wire CLOCK_n_tid0_78;


registerNbits outA (.out ({result[31], result[30], result[29], result[28], result[27], 
    result[26], result[25], result[24], result[23], result[22], result[21], result[20], 
    result[19], result[18], result[17], result[16], result[15], result[14], result[13], 
    result[12], result[11], result[10], result[9], result[8], result[7], result[6], 
    result[5], result[4], result[3], result[2], result[1], result[0]}), .en (enableOutput)
    , .inp ({\outB_reg[31] , \outB_reg[30] , \outB_reg[29] , \outB_reg[28] , \outB_reg[27] , 
    \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , \outB_reg[23] , \outB_reg[22] , 
    \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , \outB_reg[18] , \outB_reg[17] , 
    \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , \outB_reg[13] , \outB_reg[12] , 
    \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , \outB_reg[8] , \outB_reg[7] , 
    \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , 
    \outB_reg[0] }), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_6));
registerNbits__0_28 outB (.out ({result[63], result[62], result[61], result[60], 
    result[59], result[58], result[57], result[56], result[55], result[54], result[53], 
    result[52], result[51], result[50], result[49], result[48], result[47], result[46], 
    result[45], result[44], result[43], result[42], result[41], result[40], result[39], 
    result[38], result[37], result[36], result[35], result[34], result[33], result[32]})
    , .en (enableOutput), .inp ({\outA_reg[31] , \outA_reg[30] , \outA_reg[29] , 
    \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , \outA_reg[24] , 
    \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , \outA_reg[19] , 
    \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , \outA_reg[14] , 
    \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , \outA_reg[9] , 
    \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , 
    \outA_reg[2] , \outA_reg[1] , \outA_reg[0] }), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_6));
sequentialmultiplier SM (.enableOutput (enableOutput), .result ({\outA_reg[31] , 
    \outA_reg[30] , \outA_reg[29] , \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , 
    \outA_reg[25] , \outA_reg[24] , \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , 
    \outA_reg[20] , \outA_reg[19] , \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , 
    \outA_reg[15] , \outA_reg[14] , \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , 
    \outA_reg[10] , \outA_reg[9] , \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , 
    \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , \outA_reg[1] , \outA_reg[0] , \outB_reg[31] , 
    \outB_reg[30] , \outB_reg[29] , \outB_reg[28] , \outB_reg[27] , \outB_reg[26] , 
    \outB_reg[25] , \outB_reg[24] , \outB_reg[23] , \outB_reg[22] , \outB_reg[21] , 
    \outB_reg[20] , \outB_reg[19] , \outB_reg[18] , \outB_reg[17] , \outB_reg[16] , 
    \outB_reg[15] , \outB_reg[14] , \outB_reg[13] , \outB_reg[12] , \outB_reg[11] , 
    \outB_reg[10] , \outB_reg[9] , \outB_reg[8] , \outB_reg[7] , \outB_reg[6] , \outB_reg[5] , 
    \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , \outB_reg[0] }), .clk_CTS_0_PP_1 (CTS_n_tid0_6)
    , .en (en), .in1 ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , \A_reg[27] , 
    \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , \A_reg[21] , 
    \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , \A_reg[15] , 
    \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , \A_reg[9] , 
    \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , 
    \A_reg[1] , \A_reg[0] }), .in2 ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , 
    \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , 
    \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , 
    \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , 
    \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_3)
    , .clk_CTS_0_PP_15 (CLOCK_n_tid0_78), .CTSclk_CTS_0_PP_15PP_0 (clk));
registerNbits__0_25 regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , 
    \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , 
    \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , 
    \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , 
    \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .en (en), .inp ({inputB[31], inputB[30], 
    inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], inputB[24], inputB[23], 
    inputB[22], inputB[21], inputB[20], inputB[19], inputB[18], inputB[17], inputB[16], 
    inputB[15], inputB[14], inputB[13], inputB[12], inputB[11], inputB[10], inputB[9], 
    inputB[8], inputB[7], inputB[6], inputB[5], inputB[4], inputB[3], inputB[2], 
    inputB[1], inputB[0]}), .reset (reset), .clk_CTS_0_PP_11 (CLOCK_n_tid0_78));
registerNbits__0_22 regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .clk_CTS_0_PP_0 (CTS_n_tid0_3), .en (en)
    , .inp ({inputA[31], inputA[30], inputA[29], inputA[28], inputA[27], inputA[26], 
    inputA[25], inputA[24], inputA[23], inputA[22], inputA[21], inputA[20], inputA[19], 
    inputA[18], inputA[17], inputA[16], inputA[15], inputA[14], inputA[13], inputA[12], 
    inputA[11], inputA[10], inputA[9], inputA[8], inputA[7], inputA[6], inputA[5], 
    inputA[4], inputA[3], inputA[2], inputA[1], inputA[0]}), .reset (reset), .clk_CTS_0_PP_3 (CLOCK_n_tid0_78));
CLKBUF_X3 CTS_L1_tid0__c1_tid0__c14 (.Z (CLOCK_n_tid0_78), .A (clk));

endmodule //integrationMult


