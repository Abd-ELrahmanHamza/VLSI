
// 	Thu Dec 22 20:36:44 2022
//	vlsi
//	localhost.localdomain

module registerNbits (clk_CTS_1_PP_18, clk_CTS_1_PP_19, clk, reset, en, inp, out);

output [31:0] out;
output clk_CTS_1_PP_18;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_19;
wire CTS_n_tid1_5;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid1_18;
wire CTS_n_tid1_86;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (CTS_n_tid1_5), .E (n_1), .SE (1'b0 ));
INV_X4 CTS_L5_c_tid1_7 (.ZN (CTS_n_tid1_5), .A (CTS_n_tid1_18));
INV_X16 CTS_L4_c_tid1_17 (.ZN (CTS_n_tid1_18), .A (clk_CTS_1_PP_18));
INV_X8 CTS_L3_c_tid1_31 (.ZN (clk_CTS_1_PP_18), .A (CTS_n_tid1_86));
INV_X4 CTS_L2_c_tid1_32 (.ZN (CTS_n_tid1_86), .A (clk_CTS_1_PP_19));

endmodule //registerNbits

module registerNbits__6_8 (clk_CTS_1_PP_1, clk_CTS_1_PP_10, clk_CTS_1_PP_25, clk, 
    reset, en, inp, out);

output [31:0] out;
output clk_CTS_1_PP_1;
output clk_CTS_1_PP_10;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_25;
wire n_0_1;
wire slo__n10;
wire n_1;
wire CTS_n_tid1_49;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


NAND2_X1 slo__c16 (.ZN (slo__n10), .A1 (inp[31]), .A2 (n_0_1));
INV_X4 CTS_L5_c_tid1_62 (.ZN (clk_CTS_1_PP_1), .A (clk_CTS_1_PP_10));
INV_X4 i_0_1 (.ZN (n_0_1), .A (reset));
AND2_X2 i_0_32 (.ZN (n_32), .A1 (n_0_1), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_1), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_1), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_1), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_1), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_1), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_1), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_1), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_1), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_1), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_1), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_1), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_1), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_1), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_1), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_1), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_1), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_1), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_1), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_1), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_1), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_1), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_1), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_1), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_1), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_1), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_1), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_1), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_1), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_1), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_1), .A2 (inp[0]));
OR2_X4 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_49), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_49), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_49), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_49), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_49), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_49), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_49), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_49), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_49), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_49), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_49), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_49), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_49), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_49), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_49), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_49), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_49), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_49), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_49), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_49), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_49), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_49), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_49), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_49), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_49), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_49), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_49), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_49), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_49), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_49), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_49), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid1_49), .D (n_33));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n_tid1_49), .CK (clk_CTS_1_PP_1), .E (n_1), .SE (1'b0 ));
INV_X1 slo__c18 (.ZN (n_33), .A (slo__n10));
INV_X4 CTS_L4_c_tid1_70 (.ZN (clk_CTS_1_PP_10), .A (clk_CTS_1_PP_25));

endmodule //registerNbits__6_8

module registerNbits__6_5 (clk_CTS_1_PP_1, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_1;
wire n_0_0;
wire n_1;
wire CTS_n_tid0_125;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire sgo__n1;
wire sgo__n2;
wire sgo__n3;
wire sgo__n4;
wire slo__n5;
wire slo__n8;
wire slo__n11;
wire slo__n14;
wire slo__n20;
wire slo__n59;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X2 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X2 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid0_125), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (slo__n14), .CK (CTS_n_tid0_125), .D (n_3));
DFF_X2 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid0_125), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (slo__n8), .CK (CTS_n_tid0_125), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (slo__n5), .CK (CTS_n_tid0_125), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (sgo__n2), .CK (CTS_n_tid0_125), .D (n_7));
DFF_X2 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid0_125), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (sgo__n4), .CK (CTS_n_tid0_125), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (sgo__n1), .CK (CTS_n_tid0_125), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (sgo__n3), .CK (CTS_n_tid0_125), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (slo__n11), .CK (CTS_n_tid0_125), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (slo__n20), .CK (CTS_n_tid0_125), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (slo__n59), .CK (CTS_n_tid0_125), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid0_125), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid0_125), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid0_125), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid0_125), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid0_125), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid0_125), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid0_125), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid0_125), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid0_125), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid0_125), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid0_125), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid0_125), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid0_125), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid0_125), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid0_125), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid0_125), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid0_125), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid0_125), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid0_125), .D (n_33));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n_tid0_125), .CK (clk_CTS_1_PP_1), .E (n_1), .SE (1'b0 ));
BUF_X8 sgo__c1 (.Z (out[8]), .A (sgo__n1));
BUF_X8 sgo__c2 (.Z (out[5]), .A (sgo__n2));
BUF_X4 sgo__c3 (.Z (out[9]), .A (sgo__n3));
BUF_X8 sgo__c4 (.Z (out[7]), .A (sgo__n4));
BUF_X8 slo__c5 (.Z (out[4]), .A (slo__n5));
BUF_X8 slo__c8 (.Z (out[3]), .A (slo__n8));
BUF_X8 slo__c11 (.Z (out[10]), .A (slo__n11));
BUF_X4 slo__c14 (.Z (out[1]), .A (slo__n14));
BUF_X8 slo__c18 (.Z (out[11]), .A (slo__n20));
BUF_X8 slo__c37 (.Z (out[12]), .A (slo__n59));

endmodule //registerNbits__6_5

module registerNbits__6_2 (clk_CTS_1_PP_10, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_10;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_54;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire sgo__n1;
wire sgo__n2;
wire slo__n3;
wire slo__n4;
wire slo__n12;
wire slo__n15;
wire slo__n27;
wire CTS_n_tid1_62;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X2 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X2 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_54), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_54), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (sgo__n2), .CK (CTS_n_tid1_54), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (sgo__n1), .CK (CTS_n_tid1_54), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (slo__n27), .CK (CTS_n_tid1_54), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_54), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_54), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (slo__n12), .CK (CTS_n_tid1_54), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (slo__n3), .CK (CTS_n_tid1_54), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (slo__n15), .CK (CTS_n_tid1_54), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_54), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_54), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_54), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_54), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_54), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_54), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_54), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_54), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_54), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_54), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_54), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_54), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_54), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_54), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_54), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_54), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_54), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_54), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_54), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_54), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_54), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid1_54), .D (n_33));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n_tid1_54), .CK (CTS_n_tid1_62), .E (n_1), .SE (1'b0 ));
BUF_X8 sgo__c1 (.Z (out[3]), .A (sgo__n1));
BUF_X8 sgo__c2 (.Z (out[2]), .A (sgo__n2));
INV_X1 slo__c3 (.ZN (slo__n4), .A (slo__n3));
INV_X4 slo__c4 (.ZN (out[8]), .A (slo__n4));
BUF_X8 slo__c10 (.Z (out[7]), .A (slo__n12));
BUF_X4 slo__c13 (.Z (out[9]), .A (slo__n15));
BUF_X8 slo__c19 (.Z (out[4]), .A (slo__n27));
INV_X8 CTS_L5_c_tid1_45 (.ZN (CTS_n_tid1_62), .A (clk_CTS_1_PP_10));

endmodule //registerNbits__6_2

module FA (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_0;
wire n_0_1;
wire n_0_2;


INV_X1 i_0_2 (.ZN (n_0_2), .A (n_0_1));
XNOR2_X1 i_0_1 (.ZN (n_0_1), .A (x), .B (y));
INV_X2 i_0_0 (.ZN (n_0_0), .A (z));
AOI22_X2 slo__sro_c4 (.ZN (sum), .A1 (n_0_0), .A2 (n_0_1), .B1 (z), .B2 (n_0_2));

endmodule //FA

module FA__5_188 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_0;
wire n_0_1;
wire n_0_2;


NAND2_X1 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
XNOR2_X2 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X2 i_0_1 (.ZN (n_0_0), .A (y), .B1 (z), .B2 (x));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_2), .A2 (n_0_0));

endmodule //FA__5_188

module FA__5_185 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_185

module FA__5_182 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X2 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_182

module FA__5_179 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_179

module FA__5_176 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_176

module FA__5_173 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_173

module FA__5_170 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_170

module FA__5_167 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_167

module FA__5_164 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_164

module FA__5_161 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_161

module FA__5_158 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_158

module FA__5_155 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_155

module FA__5_152 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_152

module FA__5_149 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_149

module FA__5_146 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_146

module FA__5_143 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_143

module FA__5_140 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_140

module FA__5_137 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_137

module FA__5_134 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_134

module FA__5_131 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_131

module FA__5_128 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_128

module FA__5_125 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_125

module FA__5_122 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_122

module FA__5_119 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_119

module FA__5_116 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_116

module FA__5_113 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X2 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_113

module FA__5_110 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_110

module FA__5_107 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


NAND2_X1 i_0_5 (.ZN (n_0_3), .A1 (x), .A2 (y));
OR2_X1 i_0_4 (.ZN (n_0_2), .A1 (x), .A2 (y));
NAND2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (n_0_2));
NAND2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_107

module FA__5_104 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;


NOR2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (y), .B1 (z), .B2 (x));
NOR2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_104

module FA__5_101 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;


NOR2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (y), .B1 (z), .B2 (x));
NOR2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_101

module FA__5_98 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;


NOR2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (y), .B1 (z), .B2 (x));
NOR2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_98

module FA__5_95 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;


NOR2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (y), .B1 (z), .B2 (x));
NOR2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X2 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_95

module FA__5_92 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;


NOR2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (y), .B1 (z), .B2 (x));
NOR2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X2 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_92

module FA__5_89 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;


NOR2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (y), .B1 (z), .B2 (x));
NOR2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X2 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_89

module FA__5_86 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;


NOR2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
AOI21_X2 i_0_1 (.ZN (n_0_0), .A (y), .B1 (z), .B2 (x));
NOR2_X4 i_0_0 (.ZN (cout), .A1 (n_0_0), .A2 (n_0_2));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X2 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_86

module FA__5_83 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_83

module FA__5_80 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_80

module FA__5_77 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_77

module FA__5_74 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X4 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_74

module FA__5_71 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_71

module FA__5_68 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_68

module FA__5_65 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_2;
wire slo__mro_n7;


NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X2 slo__mro_c12 (.ZN (slo__mro_n7), .A (y), .B1 (z), .B2 (x));
NAND2_X4 slo__mro_c13 (.ZN (cout), .A1 (slo__mro_n7), .A2 (n_0_2));

endmodule //FA__5_65

module FA__5_62 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_62

module FA__5_59 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_59

module FA__5_56 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_56

module FA__5_53 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X4 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_53

module FA__5_50 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_2;
wire slo__mro_n7;


NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));
OAI21_X4 slo__mro_c12 (.ZN (slo__mro_n7), .A (y), .B1 (z), .B2 (x));
NAND2_X4 slo__mro_c13 (.ZN (cout), .A1 (n_0_2), .A2 (slo__mro_n7));

endmodule //FA__5_50

module FA__5_47 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_47

module FA__5_44 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_44

module FA__5_41 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_41

module FA__5_38 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_38

module FA__5_35 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire n_0_1;
wire n_0_0;
wire n_0_2;
wire n_0_3;


INV_X1 i_0_5 (.ZN (n_0_3), .A (y));
NAND2_X2 i_0_4 (.ZN (n_0_2), .A1 (z), .A2 (x));
NOR2_X2 i_0_1 (.ZN (n_0_0), .A1 (z), .A2 (x));
OAI21_X4 i_0_0 (.ZN (cout), .A (n_0_2), .B1 (n_0_0), .B2 (n_0_3));
XNOR2_X1 i_0_3 (.ZN (n_0_1), .A (z), .B (x));
XNOR2_X1 i_0_2 (.ZN (sum), .A (y), .B (n_0_1));

endmodule //FA__5_35

module FA__5_32 (x, y, z, sum, cout);

output cout;
output sum;
input x;
input y;
input z;
wire slo_n12;


AND2_X4 i_0_0 (.ZN (cout), .A1 (x), .A2 (y));
XOR2_X1 i_0_1 (.Z (sum), .A (y), .B (slo_n12));
CLKBUF_X1 slo___L1_c1_c11 (.Z (slo_n12), .A (x));

endmodule //FA__5_32

module RCA64 (A, B, cin, sum);

output [63:0] sum;
input [63:0] A;
input [63:0] B;
input cin;
wire \carry[63] ;
wire \carry[62] ;
wire \carry[61] ;
wire \carry[60] ;
wire \carry[59] ;
wire \carry[58] ;
wire \carry[57] ;
wire \carry[56] ;
wire \carry[55] ;
wire \carry[54] ;
wire \carry[53] ;
wire \carry[52] ;
wire \carry[51] ;
wire \carry[50] ;
wire \carry[49] ;
wire \carry[48] ;
wire \carry[47] ;
wire \carry[46] ;
wire \carry[45] ;
wire \carry[44] ;
wire \carry[43] ;
wire \carry[42] ;
wire \carry[41] ;
wire \carry[40] ;
wire \carry[39] ;
wire \carry[38] ;
wire \carry[37] ;
wire \carry[36] ;
wire \carry[35] ;
wire \carry[34] ;
wire \carry[33] ;
wire \carry[32] ;
wire \carry[31] ;
wire \carry[30] ;
wire \carry[29] ;
wire \carry[28] ;
wire \carry[27] ;
wire \carry[26] ;
wire \carry[25] ;
wire \carry[24] ;
wire \carry[23] ;
wire \carry[22] ;
wire \carry[21] ;
wire \carry[20] ;
wire \carry[19] ;
wire \carry[18] ;
wire \carry[17] ;
wire \carry[16] ;
wire \carry[15] ;
wire \carry[14] ;
wire \carry[13] ;
wire \carry[12] ;
wire \carry[11] ;


FA genblk1_63_Full_Adder (.sum (sum[63]), .x (A[63]), .y (B[63]), .z (\carry[63] ));
FA__5_188 genblk1_62_Full_Adder (.cout (\carry[63] ), .sum (sum[62]), .x (A[62]), .y (B[62]), .z (\carry[62] ));
FA__5_185 genblk1_61_Full_Adder (.cout (\carry[62] ), .sum (sum[61]), .x (A[61]), .y (B[61]), .z (\carry[61] ));
FA__5_182 genblk1_60_Full_Adder (.cout (\carry[61] ), .sum (sum[60]), .x (A[60]), .y (B[60])
    , .z (\carry[60] ));
FA__5_179 genblk1_59_Full_Adder (.cout (\carry[60] ), .sum (sum[59]), .x (A[59]), .y (B[59]), .z (\carry[59] ));
FA__5_176 genblk1_58_Full_Adder (.cout (\carry[59] ), .sum (sum[58]), .x (A[58]), .y (B[58]), .z (\carry[58] ));
FA__5_173 genblk1_57_Full_Adder (.cout (\carry[58] ), .sum (sum[57]), .x (A[57]), .y (B[57]), .z (\carry[57] ));
FA__5_170 genblk1_56_Full_Adder (.cout (\carry[57] ), .sum (sum[56]), .x (A[56]), .y (B[56])
    , .z (\carry[56] ));
FA__5_167 genblk1_55_Full_Adder (.cout (\carry[56] ), .sum (sum[55]), .x (A[55]), .y (B[55])
    , .z (\carry[55] ));
FA__5_164 genblk1_54_Full_Adder (.cout (\carry[55] ), .sum (sum[54]), .x (A[54]), .y (B[54]), .z (\carry[54] ));
FA__5_161 genblk1_53_Full_Adder (.cout (\carry[54] ), .sum (sum[53]), .x (A[53]), .y (B[53])
    , .z (\carry[53] ));
FA__5_158 genblk1_52_Full_Adder (.cout (\carry[53] ), .sum (sum[52]), .x (A[52]), .y (B[52]), .z (\carry[52] ));
FA__5_155 genblk1_51_Full_Adder (.cout (\carry[52] ), .sum (sum[51]), .x (A[51]), .y (B[51]), .z (\carry[51] ));
FA__5_152 genblk1_50_Full_Adder (.cout (\carry[51] ), .sum (sum[50]), .x (A[50]), .y (B[50]), .z (\carry[50] ));
FA__5_149 genblk1_49_Full_Adder (.cout (\carry[50] ), .sum (sum[49]), .x (A[49]), .y (B[49]), .z (\carry[49] ));
FA__5_146 genblk1_48_Full_Adder (.cout (\carry[49] ), .sum (sum[48]), .x (A[48]), .y (B[48]), .z (\carry[48] ));
FA__5_143 genblk1_47_Full_Adder (.cout (\carry[48] ), .sum (sum[47]), .x (A[47]), .y (B[47]), .z (\carry[47] ));
FA__5_140 genblk1_46_Full_Adder (.cout (\carry[47] ), .sum (sum[46]), .x (A[46]), .y (B[46]), .z (\carry[46] ));
FA__5_137 genblk1_45_Full_Adder (.cout (\carry[46] ), .sum (sum[45]), .x (A[45]), .y (B[45]), .z (\carry[45] ));
FA__5_134 genblk1_44_Full_Adder (.cout (\carry[45] ), .sum (sum[44]), .x (A[44]), .y (B[44]), .z (\carry[44] ));
FA__5_131 genblk1_43_Full_Adder (.cout (\carry[44] ), .sum (sum[43]), .x (A[43]), .y (B[43]), .z (\carry[43] ));
FA__5_128 genblk1_42_Full_Adder (.cout (\carry[43] ), .sum (sum[42]), .x (A[42]), .y (B[42]), .z (\carry[42] ));
FA__5_125 genblk1_41_Full_Adder (.cout (\carry[42] ), .sum (sum[41]), .x (A[41]), .y (B[41]), .z (\carry[41] ));
FA__5_122 genblk1_40_Full_Adder (.cout (\carry[41] ), .sum (sum[40]), .x (A[40]), .y (B[40]), .z (\carry[40] ));
FA__5_119 genblk1_39_Full_Adder (.cout (\carry[40] ), .sum (sum[39]), .x (A[39]), .y (B[39]), .z (\carry[39] ));
FA__5_116 genblk1_38_Full_Adder (.cout (\carry[39] ), .sum (sum[38]), .x (A[38]), .y (B[38]), .z (\carry[38] ));
FA__5_113 genblk1_37_Full_Adder (.cout (\carry[38] ), .sum (sum[37]), .x (A[37]), .y (B[37]), .z (\carry[37] ));
FA__5_110 genblk1_36_Full_Adder (.cout (\carry[37] ), .sum (sum[36]), .x (A[36]), .y (B[36]), .z (\carry[36] ));
FA__5_107 genblk1_35_Full_Adder (.cout (\carry[36] ), .sum (sum[35]), .x (A[35]), .y (B[35]), .z (\carry[35] ));
FA__5_104 genblk1_34_Full_Adder (.cout (\carry[35] ), .sum (sum[34]), .x (A[34]), .y (B[34]), .z (\carry[34] ));
FA__5_101 genblk1_33_Full_Adder (.cout (\carry[34] ), .sum (sum[33]), .x (A[33]), .y (B[33]), .z (\carry[33] ));
FA__5_98 genblk1_32_Full_Adder (.cout (\carry[33] ), .sum (sum[32]), .x (A[32]), .y (B[32]), .z (\carry[32] ));
FA__5_95 genblk1_31_Full_Adder (.cout (\carry[32] ), .sum (sum[31]), .x (A[31]), .y (B[31]), .z (\carry[31] ));
FA__5_92 genblk1_30_Full_Adder (.cout (\carry[31] ), .sum (sum[30]), .x (A[30]), .y (B[30]), .z (\carry[30] ));
FA__5_89 genblk1_29_Full_Adder (.cout (\carry[30] ), .sum (sum[29]), .x (A[29]), .y (B[29]), .z (\carry[29] ));
FA__5_86 genblk1_28_Full_Adder (.cout (\carry[29] ), .sum (sum[28]), .x (A[28]), .y (B[28]), .z (\carry[28] ));
FA__5_83 genblk1_27_Full_Adder (.cout (\carry[28] ), .sum (sum[27]), .x (A[27]), .y (B[27]), .z (\carry[27] ));
FA__5_80 genblk1_26_Full_Adder (.cout (\carry[27] ), .sum (sum[26]), .x (A[26]), .y (B[26]), .z (\carry[26] ));
FA__5_77 genblk1_25_Full_Adder (.cout (\carry[26] ), .sum (sum[25]), .x (A[25]), .y (B[25]), .z (\carry[25] ));
FA__5_74 genblk1_24_Full_Adder (.cout (\carry[25] ), .sum (sum[24]), .x (A[24]), .y (B[24]), .z (\carry[24] ));
FA__5_71 genblk1_23_Full_Adder (.cout (\carry[24] ), .sum (sum[23]), .x (A[23]), .y (B[23]), .z (\carry[23] ));
FA__5_68 genblk1_22_Full_Adder (.cout (\carry[23] ), .sum (sum[22]), .x (A[22]), .y (B[22]), .z (\carry[22] ));
FA__5_65 genblk1_21_Full_Adder (.cout (\carry[22] ), .sum (sum[21]), .x (A[21]), .y (B[21]), .z (\carry[21] ));
FA__5_62 genblk1_20_Full_Adder (.cout (\carry[21] ), .sum (sum[20]), .x (A[20]), .y (B[20]), .z (\carry[20] ));
FA__5_59 genblk1_19_Full_Adder (.cout (\carry[20] ), .sum (sum[19]), .x (A[19]), .y (B[19]), .z (\carry[19] ));
FA__5_56 genblk1_18_Full_Adder (.cout (\carry[19] ), .sum (sum[18]), .x (A[18]), .y (B[18]), .z (\carry[18] ));
FA__5_53 genblk1_17_Full_Adder (.cout (\carry[18] ), .sum (sum[17]), .x (A[17]), .y (B[17]), .z (\carry[17] ));
FA__5_50 genblk1_16_Full_Adder (.cout (\carry[17] ), .sum (sum[16]), .x (A[16]), .y (B[16]), .z (\carry[16] ));
FA__5_47 genblk1_15_Full_Adder (.cout (\carry[16] ), .sum (sum[15]), .x (A[15]), .y (B[15]), .z (\carry[15] ));
FA__5_44 genblk1_14_Full_Adder (.cout (\carry[15] ), .sum (sum[14]), .x (A[14]), .y (B[14]), .z (\carry[14] ));
FA__5_41 genblk1_13_Full_Adder (.cout (\carry[14] ), .sum (sum[13]), .x (A[13]), .y (B[13]), .z (\carry[13] ));
FA__5_38 genblk1_12_Full_Adder (.cout (\carry[13] ), .sum (sum[12]), .x (A[12]), .y (B[12]), .z (\carry[12] ));
FA__5_35 genblk1_11_Full_Adder (.cout (\carry[12] ), .sum (sum[11]), .x (A[11]), .y (B[11]), .z (\carry[11] ));
FA__5_32 genblk1_10_Full_Adder (.cout (\carry[11] ), .sum (sum[10]), .x (A[10]), .y (B[10]));

endmodule //RCA64

module CSA (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;


XOR2_X1 i_0_123 (.Z (u[63]), .A (y[63]), .B (x[63]));
XOR2_X1 i_0_122 (.Z (u[62]), .A (y[62]), .B (x[62]));
XOR2_X1 i_0_121 (.Z (u[61]), .A (y[61]), .B (x[61]));
XOR2_X1 i_0_120 (.Z (u[60]), .A (y[60]), .B (x[60]));
XOR2_X1 i_0_119 (.Z (u[59]), .A (y[59]), .B (x[59]));
XOR2_X1 i_0_118 (.Z (u[58]), .A (y[58]), .B (x[58]));
XOR2_X1 i_0_117 (.Z (u[57]), .A (y[57]), .B (x[57]));
XOR2_X1 i_0_116 (.Z (u[56]), .A (y[56]), .B (x[56]));
XOR2_X1 i_0_115 (.Z (u[55]), .A (y[55]), .B (x[55]));
XOR2_X1 i_0_114 (.Z (u[54]), .A (y[54]), .B (x[54]));
XOR2_X1 i_0_113 (.Z (u[53]), .A (y[53]), .B (x[53]));
XOR2_X1 i_0_112 (.Z (u[52]), .A (y[52]), .B (x[52]));
XOR2_X1 i_0_111 (.Z (u[51]), .A (y[51]), .B (x[51]));
XOR2_X1 i_0_110 (.Z (u[50]), .A (y[50]), .B (x[50]));
XOR2_X1 i_0_109 (.Z (u[49]), .A (y[49]), .B (x[49]));
XOR2_X1 i_0_108 (.Z (u[48]), .A (y[48]), .B (x[48]));
XOR2_X1 i_0_107 (.Z (u[47]), .A (y[47]), .B (x[47]));
XOR2_X1 i_0_106 (.Z (u[46]), .A (y[46]), .B (x[46]));
XOR2_X1 i_0_105 (.Z (u[45]), .A (y[45]), .B (x[45]));
XOR2_X1 i_0_104 (.Z (u[44]), .A (y[44]), .B (x[44]));
XOR2_X1 i_0_103 (.Z (u[43]), .A (y[43]), .B (x[43]));
XOR2_X1 i_0_102 (.Z (u[42]), .A (y[42]), .B (x[42]));
XOR2_X1 i_0_101 (.Z (u[41]), .A (y[41]), .B (x[41]));
XOR2_X1 i_0_100 (.Z (u[40]), .A (y[40]), .B (x[40]));
XOR2_X1 i_0_99 (.Z (u[39]), .A (y[39]), .B (x[39]));
XOR2_X1 i_0_98 (.Z (u[38]), .A (y[38]), .B (x[38]));
XOR2_X1 i_0_97 (.Z (u[37]), .A (y[37]), .B (x[37]));
XOR2_X1 i_0_96 (.Z (u[36]), .A (y[36]), .B (x[36]));
XOR2_X1 i_0_95 (.Z (u[35]), .A (y[35]), .B (x[35]));
XOR2_X2 i_0_94 (.Z (u[34]), .A (y[34]), .B (x[34]));
XOR2_X2 i_0_93 (.Z (u[33]), .A (y[33]), .B (x[33]));
XOR2_X2 i_0_92 (.Z (u[32]), .A (y[32]), .B (x[32]));
XNOR2_X1 i_0_91 (.ZN (n_0_2), .A (z[31]), .B (x[31]));
XNOR2_X2 i_0_90 (.ZN (u[31]), .A (y[31]), .B (n_0_2));
XOR2_X2 i_0_89 (.Z (u[30]), .A (y[30]), .B (x[30]));
XOR2_X2 i_0_88 (.Z (u[29]), .A (y[29]), .B (x[29]));
XOR2_X2 i_0_87 (.Z (u[28]), .A (y[28]), .B (x[28]));
XOR2_X2 i_0_86 (.Z (u[27]), .A (y[27]), .B (x[27]));
XOR2_X2 i_0_85 (.Z (u[26]), .A (y[26]), .B (x[26]));
XOR2_X2 i_0_84 (.Z (u[25]), .A (y[25]), .B (x[25]));
XOR2_X2 i_0_83 (.Z (u[24]), .A (y[24]), .B (x[24]));
XOR2_X2 i_0_82 (.Z (u[23]), .A (y[23]), .B (x[23]));
XOR2_X2 i_0_81 (.Z (u[22]), .A (y[22]), .B (x[22]));
XOR2_X2 i_0_80 (.Z (u[21]), .A (y[21]), .B (x[21]));
XOR2_X2 i_0_79 (.Z (u[20]), .A (y[20]), .B (x[20]));
XOR2_X2 i_0_78 (.Z (u[19]), .A (y[19]), .B (x[19]));
XOR2_X2 i_0_77 (.Z (u[18]), .A (y[18]), .B (x[18]));
XOR2_X2 i_0_76 (.Z (u[17]), .A (y[17]), .B (x[17]));
XOR2_X2 i_0_75 (.Z (u[16]), .A (y[16]), .B (x[16]));
XOR2_X2 i_0_74 (.Z (u[15]), .A (y[15]), .B (x[15]));
XOR2_X2 i_0_73 (.Z (u[14]), .A (y[14]), .B (x[14]));
XOR2_X2 i_0_72 (.Z (u[13]), .A (y[13]), .B (x[13]));
XOR2_X2 i_0_71 (.Z (u[12]), .A (y[12]), .B (x[12]));
XOR2_X2 i_0_70 (.Z (u[11]), .A (y[11]), .B (x[11]));
XOR2_X2 i_0_69 (.Z (u[10]), .A (y[10]), .B (x[10]));
XOR2_X1 i_0_68 (.Z (u[9]), .A (y[9]), .B (x[9]));
AND2_X1 i_0_61 (.ZN (v[63]), .A1 (y[62]), .A2 (x[62]));
AND2_X1 i_0_60 (.ZN (v[62]), .A1 (y[61]), .A2 (x[61]));
AND2_X1 i_0_59 (.ZN (v[61]), .A1 (y[60]), .A2 (x[60]));
AND2_X1 i_0_58 (.ZN (v[60]), .A1 (y[59]), .A2 (x[59]));
AND2_X1 i_0_57 (.ZN (v[59]), .A1 (y[58]), .A2 (x[58]));
AND2_X1 i_0_56 (.ZN (v[58]), .A1 (y[57]), .A2 (x[57]));
AND2_X1 i_0_55 (.ZN (v[57]), .A1 (y[56]), .A2 (x[56]));
AND2_X1 i_0_54 (.ZN (v[56]), .A1 (y[55]), .A2 (x[55]));
AND2_X1 i_0_53 (.ZN (v[55]), .A1 (y[54]), .A2 (x[54]));
AND2_X1 i_0_52 (.ZN (v[54]), .A1 (y[53]), .A2 (x[53]));
AND2_X1 i_0_51 (.ZN (v[53]), .A1 (y[52]), .A2 (x[52]));
AND2_X1 i_0_50 (.ZN (v[52]), .A1 (y[51]), .A2 (x[51]));
AND2_X1 i_0_49 (.ZN (v[51]), .A1 (y[50]), .A2 (x[50]));
AND2_X1 i_0_48 (.ZN (v[50]), .A1 (y[49]), .A2 (x[49]));
AND2_X1 i_0_47 (.ZN (v[49]), .A1 (y[48]), .A2 (x[48]));
AND2_X1 i_0_46 (.ZN (v[48]), .A1 (y[47]), .A2 (x[47]));
AND2_X1 i_0_45 (.ZN (v[47]), .A1 (y[46]), .A2 (x[46]));
AND2_X1 i_0_44 (.ZN (v[46]), .A1 (y[45]), .A2 (x[45]));
AND2_X1 i_0_43 (.ZN (v[45]), .A1 (y[44]), .A2 (x[44]));
AND2_X1 i_0_42 (.ZN (v[44]), .A1 (y[43]), .A2 (x[43]));
AND2_X1 i_0_41 (.ZN (v[43]), .A1 (y[42]), .A2 (x[42]));
AND2_X1 i_0_40 (.ZN (v[42]), .A1 (y[41]), .A2 (x[41]));
AND2_X1 i_0_39 (.ZN (v[41]), .A1 (y[40]), .A2 (x[40]));
AND2_X1 i_0_38 (.ZN (v[40]), .A1 (y[39]), .A2 (x[39]));
AND2_X1 i_0_37 (.ZN (v[39]), .A1 (y[38]), .A2 (x[38]));
AND2_X1 i_0_36 (.ZN (v[38]), .A1 (y[37]), .A2 (x[37]));
AND2_X1 i_0_35 (.ZN (v[37]), .A1 (y[36]), .A2 (x[36]));
AND2_X1 i_0_34 (.ZN (v[36]), .A1 (y[35]), .A2 (x[35]));
AND2_X1 i_0_33 (.ZN (v[35]), .A1 (y[34]), .A2 (x[34]));
AND2_X1 i_0_32 (.ZN (v[34]), .A1 (y[33]), .A2 (x[33]));
AND2_X1 i_0_31 (.ZN (v[33]), .A1 (y[32]), .A2 (x[32]));
NAND2_X1 i_0_30 (.ZN (n_0_1), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_29 (.ZN (n_0_0), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_28 (.ZN (v[32]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_27 (.ZN (v[31]), .A1 (y[30]), .A2 (x[30]));
AND2_X1 i_0_26 (.ZN (v[30]), .A1 (y[29]), .A2 (x[29]));
AND2_X1 i_0_25 (.ZN (v[29]), .A1 (y[28]), .A2 (x[28]));
AND2_X1 i_0_24 (.ZN (v[28]), .A1 (y[27]), .A2 (x[27]));
AND2_X1 i_0_23 (.ZN (v[27]), .A1 (y[26]), .A2 (x[26]));
AND2_X1 i_0_22 (.ZN (v[26]), .A1 (y[25]), .A2 (x[25]));
AND2_X1 i_0_21 (.ZN (v[25]), .A1 (y[24]), .A2 (x[24]));
AND2_X1 i_0_20 (.ZN (v[24]), .A1 (y[23]), .A2 (x[23]));
AND2_X1 i_0_19 (.ZN (v[23]), .A1 (y[22]), .A2 (x[22]));
AND2_X1 i_0_18 (.ZN (v[22]), .A1 (y[21]), .A2 (x[21]));
AND2_X1 i_0_17 (.ZN (v[21]), .A1 (y[20]), .A2 (x[20]));
AND2_X1 i_0_16 (.ZN (v[20]), .A1 (y[19]), .A2 (x[19]));
AND2_X1 i_0_15 (.ZN (v[19]), .A1 (y[18]), .A2 (x[18]));
AND2_X1 i_0_14 (.ZN (v[18]), .A1 (y[17]), .A2 (x[17]));
AND2_X1 i_0_13 (.ZN (v[17]), .A1 (y[16]), .A2 (x[16]));
AND2_X1 i_0_12 (.ZN (v[16]), .A1 (y[15]), .A2 (x[15]));
AND2_X1 i_0_11 (.ZN (v[15]), .A1 (y[14]), .A2 (x[14]));
AND2_X1 i_0_10 (.ZN (v[14]), .A1 (y[13]), .A2 (x[13]));
AND2_X1 i_0_9 (.ZN (v[13]), .A1 (y[12]), .A2 (x[12]));
AND2_X1 i_0_8 (.ZN (v[12]), .A1 (y[11]), .A2 (x[11]));
AND2_X1 i_0_7 (.ZN (v[11]), .A1 (y[10]), .A2 (x[10]));
AND2_X4 i_0_6 (.ZN (v[10]), .A1 (y[9]), .A2 (x[9]));

endmodule //CSA

module CSA__5_212 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;


XNOR2_X1 i_0_219 (.ZN (n_0_96), .A (z[63]), .B (x[63]));
XNOR2_X1 i_0_218 (.ZN (u[63]), .A (y[63]), .B (n_0_96));
XNOR2_X1 i_0_217 (.ZN (n_0_95), .A (z[62]), .B (x[62]));
XNOR2_X1 i_0_216 (.ZN (u[62]), .A (y[62]), .B (n_0_95));
XNOR2_X1 i_0_215 (.ZN (n_0_94), .A (z[61]), .B (x[61]));
XNOR2_X1 i_0_214 (.ZN (u[61]), .A (y[61]), .B (n_0_94));
XNOR2_X1 i_0_213 (.ZN (n_0_93), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_212 (.ZN (u[60]), .A (y[60]), .B (n_0_93));
XNOR2_X1 i_0_211 (.ZN (n_0_92), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_210 (.ZN (u[59]), .A (y[59]), .B (n_0_92));
XNOR2_X1 i_0_209 (.ZN (n_0_91), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_208 (.ZN (u[58]), .A (y[58]), .B (n_0_91));
XNOR2_X1 i_0_207 (.ZN (n_0_90), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_206 (.ZN (u[57]), .A (y[57]), .B (n_0_90));
XNOR2_X1 i_0_205 (.ZN (n_0_89), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_204 (.ZN (u[56]), .A (y[56]), .B (n_0_89));
XNOR2_X1 i_0_203 (.ZN (n_0_88), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_202 (.ZN (u[55]), .A (y[55]), .B (n_0_88));
XNOR2_X1 i_0_201 (.ZN (n_0_87), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_200 (.ZN (u[54]), .A (y[54]), .B (n_0_87));
XNOR2_X1 i_0_199 (.ZN (n_0_86), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_198 (.ZN (u[53]), .A (y[53]), .B (n_0_86));
XNOR2_X1 i_0_197 (.ZN (n_0_85), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_196 (.ZN (u[52]), .A (y[52]), .B (n_0_85));
XNOR2_X1 i_0_195 (.ZN (n_0_84), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_194 (.ZN (u[51]), .A (y[51]), .B (n_0_84));
XNOR2_X1 i_0_193 (.ZN (n_0_83), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_192 (.ZN (u[50]), .A (y[50]), .B (n_0_83));
XNOR2_X1 i_0_191 (.ZN (n_0_82), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_190 (.ZN (u[49]), .A (y[49]), .B (n_0_82));
XNOR2_X1 i_0_189 (.ZN (n_0_81), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_188 (.ZN (u[48]), .A (y[48]), .B (n_0_81));
XNOR2_X1 i_0_187 (.ZN (n_0_80), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_186 (.ZN (u[47]), .A (y[47]), .B (n_0_80));
XNOR2_X1 i_0_185 (.ZN (n_0_79), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_184 (.ZN (u[46]), .A (y[46]), .B (n_0_79));
XNOR2_X1 i_0_183 (.ZN (n_0_78), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_182 (.ZN (u[45]), .A (y[45]), .B (n_0_78));
XNOR2_X1 i_0_181 (.ZN (n_0_77), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_180 (.ZN (u[44]), .A (y[44]), .B (n_0_77));
XNOR2_X1 i_0_179 (.ZN (n_0_76), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_178 (.ZN (u[43]), .A (y[43]), .B (n_0_76));
XNOR2_X1 i_0_177 (.ZN (n_0_75), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_176 (.ZN (u[42]), .A (y[42]), .B (n_0_75));
XNOR2_X1 i_0_175 (.ZN (n_0_74), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_174 (.ZN (u[41]), .A (y[41]), .B (n_0_74));
XNOR2_X1 i_0_173 (.ZN (n_0_73), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_172 (.ZN (u[40]), .A (y[40]), .B (n_0_73));
XNOR2_X1 i_0_171 (.ZN (n_0_72), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_170 (.ZN (u[39]), .A (y[39]), .B (n_0_72));
XNOR2_X1 i_0_169 (.ZN (n_0_71), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_168 (.ZN (u[38]), .A (y[38]), .B (n_0_71));
XNOR2_X1 i_0_167 (.ZN (n_0_70), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_166 (.ZN (u[37]), .A (y[37]), .B (n_0_70));
XNOR2_X1 i_0_165 (.ZN (n_0_69), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_164 (.ZN (u[36]), .A (y[36]), .B (n_0_69));
XNOR2_X1 i_0_163 (.ZN (n_0_68), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_162 (.ZN (u[35]), .A (y[35]), .B (n_0_68));
XNOR2_X1 i_0_161 (.ZN (n_0_67), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_160 (.ZN (u[34]), .A (y[34]), .B (n_0_67));
XNOR2_X1 i_0_159 (.ZN (n_0_66), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_158 (.ZN (u[33]), .A (y[33]), .B (n_0_66));
XNOR2_X1 i_0_157 (.ZN (n_0_65), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_156 (.ZN (u[32]), .A (y[32]), .B (n_0_65));
XNOR2_X1 i_0_155 (.ZN (n_0_64), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_154 (.ZN (u[31]), .A (y[31]), .B (n_0_64));
XOR2_X1 i_0_153 (.Z (u[30]), .A (y[30]), .B (x[30]));
XOR2_X1 i_0_152 (.Z (u[29]), .A (y[29]), .B (x[29]));
XOR2_X1 i_0_151 (.Z (u[28]), .A (y[28]), .B (x[28]));
XOR2_X1 i_0_150 (.Z (u[27]), .A (y[27]), .B (x[27]));
XOR2_X1 i_0_149 (.Z (u[26]), .A (y[26]), .B (x[26]));
XOR2_X1 i_0_148 (.Z (u[25]), .A (y[25]), .B (x[25]));
XOR2_X1 i_0_147 (.Z (u[24]), .A (y[24]), .B (x[24]));
XOR2_X1 i_0_146 (.Z (u[23]), .A (y[23]), .B (x[23]));
XOR2_X1 i_0_145 (.Z (u[22]), .A (y[22]), .B (x[22]));
XOR2_X1 i_0_144 (.Z (u[21]), .A (y[21]), .B (x[21]));
XOR2_X1 i_0_143 (.Z (u[20]), .A (y[20]), .B (x[20]));
XOR2_X1 i_0_142 (.Z (u[19]), .A (y[19]), .B (x[19]));
XOR2_X1 i_0_141 (.Z (u[18]), .A (y[18]), .B (x[18]));
XOR2_X1 i_0_140 (.Z (u[17]), .A (y[17]), .B (x[17]));
XOR2_X1 i_0_139 (.Z (u[16]), .A (y[16]), .B (x[16]));
XOR2_X2 i_0_138 (.Z (u[15]), .A (y[15]), .B (x[15]));
XOR2_X2 i_0_137 (.Z (u[14]), .A (y[14]), .B (x[14]));
XOR2_X2 i_0_136 (.Z (u[13]), .A (y[13]), .B (x[13]));
XOR2_X2 i_0_135 (.Z (u[12]), .A (y[12]), .B (x[12]));
XOR2_X2 i_0_134 (.Z (u[11]), .A (y[11]), .B (x[11]));
XOR2_X2 i_0_133 (.Z (u[10]), .A (y[10]), .B (x[10]));
XOR2_X2 i_0_132 (.Z (u[9]), .A (y[9]), .B (x[9]));
XOR2_X1 i_0_131 (.Z (u[8]), .A (y[8]), .B (x[8]));
NAND2_X1 i_0_124 (.ZN (n_0_63), .A1 (z[62]), .A2 (x[62]));
OAI21_X1 i_0_123 (.ZN (n_0_62), .A (y[62]), .B1 (z[62]), .B2 (x[62]));
NAND2_X1 i_0_122 (.ZN (v[63]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_121 (.ZN (n_0_61), .A1 (z[61]), .A2 (x[61]));
OAI21_X1 i_0_120 (.ZN (n_0_60), .A (y[61]), .B1 (z[61]), .B2 (x[61]));
NAND2_X1 i_0_119 (.ZN (v[62]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_118 (.ZN (n_0_59), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_117 (.ZN (n_0_58), .A (y[60]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_116 (.ZN (v[61]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_115 (.ZN (n_0_57), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_114 (.ZN (n_0_56), .A (y[59]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_113 (.ZN (v[60]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_112 (.ZN (n_0_55), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_111 (.ZN (n_0_54), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_110 (.ZN (v[59]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_109 (.ZN (n_0_53), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_108 (.ZN (n_0_52), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_107 (.ZN (v[58]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_106 (.ZN (n_0_51), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_105 (.ZN (n_0_50), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_104 (.ZN (v[57]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_103 (.ZN (n_0_49), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_102 (.ZN (n_0_48), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_101 (.ZN (v[56]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_100 (.ZN (n_0_47), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_99 (.ZN (n_0_46), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_98 (.ZN (v[55]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_97 (.ZN (n_0_45), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_96 (.ZN (n_0_44), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_95 (.ZN (v[54]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_94 (.ZN (n_0_43), .A1 (y[52]), .A2 (x[52]));
OAI21_X1 i_0_93 (.ZN (n_0_42), .A (z[52]), .B1 (x[52]), .B2 (y[52]));
NAND2_X1 i_0_92 (.ZN (v[53]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_91 (.ZN (n_0_41), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_90 (.ZN (n_0_40), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_89 (.ZN (v[52]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_88 (.ZN (n_0_39), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_87 (.ZN (n_0_38), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_86 (.ZN (v[51]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_85 (.ZN (n_0_37), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_84 (.ZN (n_0_36), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_83 (.ZN (v[50]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_82 (.ZN (n_0_35), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_81 (.ZN (n_0_34), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_80 (.ZN (v[49]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_79 (.ZN (n_0_33), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_78 (.ZN (n_0_32), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_77 (.ZN (v[48]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_76 (.ZN (n_0_31), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_75 (.ZN (n_0_30), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_74 (.ZN (v[47]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_73 (.ZN (n_0_29), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_72 (.ZN (n_0_28), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_71 (.ZN (v[46]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_70 (.ZN (n_0_27), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_69 (.ZN (n_0_26), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_68 (.ZN (v[45]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_67 (.ZN (n_0_25), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_66 (.ZN (n_0_24), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_65 (.ZN (v[44]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_64 (.ZN (n_0_23), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_63 (.ZN (n_0_22), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_62 (.ZN (v[43]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_61 (.ZN (n_0_21), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_60 (.ZN (n_0_20), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_59 (.ZN (v[42]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_58 (.ZN (n_0_19), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_57 (.ZN (n_0_18), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_56 (.ZN (v[41]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_55 (.ZN (n_0_17), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_54 (.ZN (n_0_16), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_53 (.ZN (v[40]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_52 (.ZN (n_0_15), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_51 (.ZN (n_0_14), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_50 (.ZN (v[39]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_49 (.ZN (n_0_13), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_48 (.ZN (n_0_12), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_47 (.ZN (v[38]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_46 (.ZN (n_0_11), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_45 (.ZN (n_0_10), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_44 (.ZN (v[37]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_43 (.ZN (n_0_9), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_42 (.ZN (n_0_8), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_41 (.ZN (v[36]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_40 (.ZN (n_0_7), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_39 (.ZN (n_0_6), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_38 (.ZN (v[35]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_37 (.ZN (n_0_5), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_36 (.ZN (n_0_4), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_35 (.ZN (v[34]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_34 (.ZN (n_0_3), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_33 (.ZN (n_0_2), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_32 (.ZN (v[33]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_31 (.ZN (n_0_1), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_30 (.ZN (n_0_0), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_29 (.ZN (v[32]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_28 (.ZN (v[31]), .A1 (y[30]), .A2 (x[30]));
AND2_X1 i_0_27 (.ZN (v[30]), .A1 (y[29]), .A2 (x[29]));
AND2_X1 i_0_26 (.ZN (v[29]), .A1 (y[28]), .A2 (x[28]));
AND2_X1 i_0_25 (.ZN (v[28]), .A1 (y[27]), .A2 (x[27]));
AND2_X1 i_0_24 (.ZN (v[27]), .A1 (y[26]), .A2 (x[26]));
AND2_X1 i_0_23 (.ZN (v[26]), .A1 (y[25]), .A2 (x[25]));
AND2_X1 i_0_22 (.ZN (v[25]), .A1 (y[24]), .A2 (x[24]));
AND2_X1 i_0_21 (.ZN (v[24]), .A1 (y[23]), .A2 (x[23]));
AND2_X1 i_0_20 (.ZN (v[23]), .A1 (y[22]), .A2 (x[22]));
AND2_X1 i_0_19 (.ZN (v[22]), .A1 (y[21]), .A2 (x[21]));
AND2_X1 i_0_18 (.ZN (v[21]), .A1 (y[20]), .A2 (x[20]));
AND2_X1 i_0_17 (.ZN (v[20]), .A1 (y[19]), .A2 (x[19]));
AND2_X1 i_0_16 (.ZN (v[19]), .A1 (y[18]), .A2 (x[18]));
AND2_X1 i_0_15 (.ZN (v[18]), .A1 (y[17]), .A2 (x[17]));
AND2_X1 i_0_14 (.ZN (v[17]), .A1 (y[16]), .A2 (x[16]));
AND2_X1 i_0_13 (.ZN (v[16]), .A1 (y[15]), .A2 (x[15]));
AND2_X1 i_0_12 (.ZN (v[15]), .A1 (y[14]), .A2 (x[14]));
AND2_X1 i_0_11 (.ZN (v[14]), .A1 (y[13]), .A2 (x[13]));
AND2_X1 i_0_10 (.ZN (v[13]), .A1 (y[12]), .A2 (x[12]));
AND2_X1 i_0_9 (.ZN (v[12]), .A1 (y[11]), .A2 (x[11]));
AND2_X1 i_0_8 (.ZN (v[11]), .A1 (y[10]), .A2 (x[10]));
AND2_X2 i_0_7 (.ZN (v[10]), .A1 (y[9]), .A2 (x[9]));
AND2_X4 i_0_6 (.ZN (v[9]), .A1 (y[8]), .A2 (x[8]));

endmodule //CSA__5_212

module CSA__5_209 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire slo_n27;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;


XOR2_X2 i_0_0 (.Z (u[10]), .A (y[10]), .B (x[10]));
XNOR2_X1 i_0_246 (.ZN (n_0_123), .A (z[63]), .B (x[63]));
XNOR2_X1 i_0_245 (.ZN (u[63]), .A (y[63]), .B (n_0_123));
XNOR2_X1 i_0_244 (.ZN (n_0_122), .A (z[62]), .B (x[62]));
XNOR2_X1 i_0_243 (.ZN (u[62]), .A (y[62]), .B (n_0_122));
XNOR2_X1 i_0_242 (.ZN (n_0_121), .A (z[61]), .B (x[61]));
XNOR2_X1 i_0_241 (.ZN (u[61]), .A (y[61]), .B (n_0_121));
XNOR2_X1 i_0_240 (.ZN (n_0_120), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_239 (.ZN (u[60]), .A (y[60]), .B (n_0_120));
XNOR2_X1 i_0_238 (.ZN (n_0_119), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_237 (.ZN (u[59]), .A (y[59]), .B (n_0_119));
XNOR2_X1 i_0_236 (.ZN (n_0_118), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_235 (.ZN (u[58]), .A (y[58]), .B (n_0_118));
XNOR2_X1 i_0_234 (.ZN (n_0_117), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_233 (.ZN (u[57]), .A (y[57]), .B (n_0_117));
XNOR2_X1 i_0_232 (.ZN (n_0_116), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_231 (.ZN (u[56]), .A (y[56]), .B (n_0_116));
XNOR2_X1 i_0_230 (.ZN (n_0_115), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_229 (.ZN (u[55]), .A (y[55]), .B (n_0_115));
XNOR2_X1 i_0_228 (.ZN (n_0_114), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_227 (.ZN (u[54]), .A (y[54]), .B (n_0_114));
XNOR2_X1 i_0_226 (.ZN (n_0_113), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_225 (.ZN (u[53]), .A (y[53]), .B (n_0_113));
XNOR2_X1 i_0_224 (.ZN (n_0_112), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_223 (.ZN (u[52]), .A (y[52]), .B (n_0_112));
XNOR2_X1 i_0_222 (.ZN (n_0_111), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_221 (.ZN (u[51]), .A (y[51]), .B (n_0_111));
XNOR2_X1 i_0_220 (.ZN (n_0_110), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_219 (.ZN (u[50]), .A (y[50]), .B (n_0_110));
XNOR2_X1 i_0_218 (.ZN (n_0_109), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_217 (.ZN (u[49]), .A (y[49]), .B (n_0_109));
XNOR2_X1 i_0_216 (.ZN (n_0_108), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_215 (.ZN (u[48]), .A (y[48]), .B (n_0_108));
XNOR2_X1 i_0_214 (.ZN (n_0_107), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_213 (.ZN (u[47]), .A (y[47]), .B (n_0_107));
XNOR2_X1 i_0_212 (.ZN (n_0_106), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_211 (.ZN (u[46]), .A (y[46]), .B (n_0_106));
XNOR2_X1 i_0_210 (.ZN (n_0_105), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_209 (.ZN (u[45]), .A (y[45]), .B (n_0_105));
XNOR2_X1 i_0_208 (.ZN (n_0_104), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_207 (.ZN (u[44]), .A (y[44]), .B (n_0_104));
XNOR2_X1 i_0_206 (.ZN (n_0_103), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_205 (.ZN (u[43]), .A (y[43]), .B (n_0_103));
XNOR2_X1 i_0_204 (.ZN (n_0_102), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_203 (.ZN (u[42]), .A (y[42]), .B (n_0_102));
XNOR2_X1 i_0_202 (.ZN (n_0_101), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_201 (.ZN (u[41]), .A (y[41]), .B (n_0_101));
XNOR2_X1 i_0_200 (.ZN (n_0_100), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_199 (.ZN (u[40]), .A (y[40]), .B (n_0_100));
XNOR2_X1 i_0_198 (.ZN (n_0_99), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_197 (.ZN (u[39]), .A (y[39]), .B (n_0_99));
XNOR2_X1 i_0_196 (.ZN (n_0_98), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_195 (.ZN (u[38]), .A (y[38]), .B (n_0_98));
XNOR2_X1 i_0_194 (.ZN (n_0_97), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_193 (.ZN (u[37]), .A (y[37]), .B (n_0_97));
XNOR2_X1 i_0_192 (.ZN (n_0_96), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_191 (.ZN (u[36]), .A (y[36]), .B (n_0_96));
XNOR2_X1 i_0_190 (.ZN (n_0_95), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_189 (.ZN (u[35]), .A (y[35]), .B (n_0_95));
XNOR2_X1 i_0_188 (.ZN (n_0_94), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_187 (.ZN (u[34]), .A (y[34]), .B (n_0_94));
XNOR2_X1 i_0_186 (.ZN (n_0_93), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_185 (.ZN (u[33]), .A (y[33]), .B (n_0_93));
XNOR2_X1 i_0_184 (.ZN (n_0_92), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_183 (.ZN (u[32]), .A (y[32]), .B (n_0_92));
XNOR2_X1 i_0_182 (.ZN (n_0_91), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_181 (.ZN (u[31]), .A (y[31]), .B (n_0_91));
XNOR2_X1 i_0_180 (.ZN (n_0_90), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_179 (.ZN (u[30]), .A (y[30]), .B (n_0_90));
XNOR2_X1 i_0_178 (.ZN (n_0_89), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_177 (.ZN (u[29]), .A (y[29]), .B (n_0_89));
XNOR2_X1 i_0_176 (.ZN (n_0_88), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_175 (.ZN (u[28]), .A (y[28]), .B (n_0_88));
XNOR2_X1 i_0_174 (.ZN (n_0_87), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_173 (.ZN (u[27]), .A (y[27]), .B (n_0_87));
XNOR2_X1 i_0_172 (.ZN (n_0_86), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_171 (.ZN (u[26]), .A (y[26]), .B (n_0_86));
XNOR2_X1 i_0_170 (.ZN (n_0_85), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_169 (.ZN (u[25]), .A (y[25]), .B (n_0_85));
XNOR2_X1 i_0_168 (.ZN (n_0_84), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_167 (.ZN (u[24]), .A (y[24]), .B (n_0_84));
XNOR2_X1 i_0_166 (.ZN (n_0_83), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_165 (.ZN (u[23]), .A (y[23]), .B (n_0_83));
XNOR2_X1 i_0_164 (.ZN (n_0_82), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_163 (.ZN (u[22]), .A (y[22]), .B (n_0_82));
XOR2_X1 i_0_162 (.Z (u[21]), .A (y[21]), .B (x[21]));
XOR2_X1 i_0_161 (.Z (u[20]), .A (y[20]), .B (x[20]));
XOR2_X1 i_0_160 (.Z (u[19]), .A (y[19]), .B (x[19]));
XOR2_X1 i_0_159 (.Z (u[18]), .A (y[18]), .B (x[18]));
XOR2_X1 i_0_158 (.Z (u[17]), .A (y[17]), .B (x[17]));
XOR2_X1 i_0_157 (.Z (u[16]), .A (y[16]), .B (x[16]));
XOR2_X2 i_0_156 (.Z (u[15]), .A (y[15]), .B (x[15]));
XOR2_X2 i_0_155 (.Z (u[14]), .A (y[14]), .B (x[14]));
XOR2_X2 i_0_154 (.Z (u[13]), .A (y[13]), .B (x[13]));
XOR2_X2 i_0_153 (.Z (u[12]), .A (y[12]), .B (x[12]));
XOR2_X2 i_0_152 (.Z (u[11]), .A (y[11]), .B (x[11]));
XOR2_X2 i_0_150 (.Z (u[9]), .A (y[9]), .B (x[9]));
XOR2_X2 i_0_149 (.Z (u[8]), .A (y[8]), .B (x[8]));
XOR2_X1 i_0_148 (.Z (u[7]), .A (y[7]), .B (x[7]));
NAND2_X1 i_0_142 (.ZN (n_0_81), .A1 (z[62]), .A2 (x[62]));
OAI21_X1 i_0_141 (.ZN (n_0_80), .A (y[62]), .B1 (z[62]), .B2 (x[62]));
NAND2_X1 i_0_140 (.ZN (v[63]), .A1 (n_0_81), .A2 (n_0_80));
NAND2_X1 i_0_139 (.ZN (n_0_79), .A1 (z[61]), .A2 (x[61]));
OAI21_X1 i_0_138 (.ZN (n_0_78), .A (y[61]), .B1 (z[61]), .B2 (x[61]));
NAND2_X1 i_0_137 (.ZN (v[62]), .A1 (n_0_79), .A2 (n_0_78));
NAND2_X1 i_0_136 (.ZN (n_0_77), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_135 (.ZN (n_0_76), .A (y[60]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_134 (.ZN (v[61]), .A1 (n_0_77), .A2 (n_0_76));
NAND2_X1 i_0_133 (.ZN (n_0_75), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_132 (.ZN (n_0_74), .A (y[59]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_131 (.ZN (v[60]), .A1 (n_0_75), .A2 (n_0_74));
NAND2_X1 i_0_130 (.ZN (n_0_73), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_129 (.ZN (n_0_72), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_128 (.ZN (v[59]), .A1 (n_0_73), .A2 (n_0_72));
NAND2_X1 i_0_127 (.ZN (n_0_71), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_126 (.ZN (n_0_70), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_125 (.ZN (v[58]), .A1 (n_0_71), .A2 (n_0_70));
NAND2_X1 i_0_124 (.ZN (n_0_69), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_123 (.ZN (n_0_68), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_122 (.ZN (v[57]), .A1 (n_0_69), .A2 (n_0_68));
NAND2_X1 i_0_121 (.ZN (n_0_67), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_120 (.ZN (n_0_66), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_119 (.ZN (v[56]), .A1 (n_0_67), .A2 (n_0_66));
NAND2_X1 i_0_118 (.ZN (n_0_65), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_117 (.ZN (n_0_64), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_116 (.ZN (v[55]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_115 (.ZN (n_0_63), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_114 (.ZN (n_0_62), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_113 (.ZN (v[54]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_112 (.ZN (n_0_61), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_111 (.ZN (n_0_60), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_110 (.ZN (v[53]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_109 (.ZN (n_0_59), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_108 (.ZN (n_0_58), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_107 (.ZN (v[52]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_106 (.ZN (n_0_57), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_105 (.ZN (n_0_56), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_104 (.ZN (v[51]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_103 (.ZN (n_0_55), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_102 (.ZN (n_0_54), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_101 (.ZN (v[50]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_100 (.ZN (n_0_53), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_99 (.ZN (n_0_52), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_98 (.ZN (v[49]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_97 (.ZN (n_0_51), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_96 (.ZN (n_0_50), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_95 (.ZN (v[48]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_94 (.ZN (n_0_49), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_93 (.ZN (n_0_48), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_92 (.ZN (v[47]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_91 (.ZN (n_0_47), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_90 (.ZN (n_0_46), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_89 (.ZN (v[46]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_88 (.ZN (n_0_45), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_87 (.ZN (n_0_44), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_86 (.ZN (v[45]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_85 (.ZN (n_0_43), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_84 (.ZN (n_0_42), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_83 (.ZN (v[44]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_82 (.ZN (n_0_41), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_81 (.ZN (n_0_40), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_80 (.ZN (v[43]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_79 (.ZN (n_0_39), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_78 (.ZN (n_0_38), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_77 (.ZN (v[42]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_76 (.ZN (n_0_37), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_75 (.ZN (n_0_36), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_74 (.ZN (v[41]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_73 (.ZN (n_0_35), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_72 (.ZN (n_0_34), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_71 (.ZN (v[40]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_70 (.ZN (n_0_33), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_69 (.ZN (n_0_32), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_68 (.ZN (v[39]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_67 (.ZN (n_0_31), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_66 (.ZN (n_0_30), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_65 (.ZN (v[38]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_64 (.ZN (n_0_29), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_63 (.ZN (n_0_28), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_62 (.ZN (v[37]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_61 (.ZN (n_0_27), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_60 (.ZN (n_0_26), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_59 (.ZN (v[36]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_58 (.ZN (n_0_25), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_57 (.ZN (n_0_24), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_56 (.ZN (v[35]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_55 (.ZN (n_0_23), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_54 (.ZN (n_0_22), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_53 (.ZN (v[34]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_52 (.ZN (n_0_21), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_51 (.ZN (n_0_20), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_50 (.ZN (v[33]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_49 (.ZN (n_0_19), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_48 (.ZN (n_0_18), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_47 (.ZN (v[32]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_46 (.ZN (n_0_17), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_45 (.ZN (n_0_16), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_44 (.ZN (v[31]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_43 (.ZN (n_0_15), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_42 (.ZN (n_0_14), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_41 (.ZN (v[30]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_40 (.ZN (n_0_13), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_39 (.ZN (n_0_12), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_38 (.ZN (v[29]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_37 (.ZN (n_0_11), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_36 (.ZN (n_0_10), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_35 (.ZN (v[28]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_34 (.ZN (n_0_9), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_33 (.ZN (n_0_8), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_32 (.ZN (v[27]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_31 (.ZN (n_0_7), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_30 (.ZN (n_0_6), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_29 (.ZN (v[26]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_28 (.ZN (n_0_5), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_27 (.ZN (n_0_4), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_26 (.ZN (v[25]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_25 (.ZN (n_0_3), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_24 (.ZN (n_0_2), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_23 (.ZN (v[24]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_22 (.ZN (n_0_1), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_21 (.ZN (n_0_0), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_20 (.ZN (v[23]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_19 (.ZN (v[22]), .A1 (y[21]), .A2 (x[21]));
AND2_X1 i_0_18 (.ZN (v[21]), .A1 (y[20]), .A2 (x[20]));
AND2_X1 i_0_17 (.ZN (v[20]), .A1 (y[19]), .A2 (x[19]));
AND2_X1 i_0_16 (.ZN (v[19]), .A1 (y[18]), .A2 (x[18]));
AND2_X1 i_0_15 (.ZN (v[18]), .A1 (y[17]), .A2 (x[17]));
AND2_X1 i_0_14 (.ZN (v[17]), .A1 (y[16]), .A2 (x[16]));
AND2_X1 i_0_13 (.ZN (v[16]), .A1 (y[15]), .A2 (x[15]));
AND2_X1 i_0_12 (.ZN (v[15]), .A1 (y[14]), .A2 (x[14]));
AND2_X1 i_0_11 (.ZN (v[14]), .A1 (y[13]), .A2 (x[13]));
AND2_X1 i_0_10 (.ZN (v[13]), .A1 (y[12]), .A2 (x[12]));
AND2_X2 i_0_9 (.ZN (v[12]), .A1 (slo_n27), .A2 (x[11]));
AND2_X1 i_0_8 (.ZN (v[11]), .A1 (y[10]), .A2 (x[10]));
AND2_X2 i_0_7 (.ZN (v[10]), .A1 (y[9]), .A2 (x[9]));
AND2_X2 i_0_6 (.ZN (v[9]), .A1 (y[8]), .A2 (x[8]));
AND2_X4 i_0_5 (.ZN (v[8]), .A1 (y[7]), .A2 (x[7]));
CLKBUF_X1 slo___L1_c1_c29 (.Z (slo_n27), .A (y[11]));

endmodule //CSA__5_209

module CSA__5_206 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire slo__mro_n9;


XOR2_X2 i_0_0 (.Z (u[10]), .A (x[10]), .B (y[10]));
XNOR2_X1 i_0_269 (.ZN (n_0_144), .A (z[63]), .B (x[63]));
XNOR2_X1 i_0_268 (.ZN (u[63]), .A (y[63]), .B (n_0_144));
XNOR2_X1 i_0_267 (.ZN (n_0_143), .A (z[62]), .B (x[62]));
XNOR2_X1 i_0_266 (.ZN (u[62]), .A (y[62]), .B (n_0_143));
XNOR2_X1 i_0_265 (.ZN (n_0_142), .A (z[61]), .B (x[61]));
XNOR2_X1 i_0_264 (.ZN (u[61]), .A (y[61]), .B (n_0_142));
XNOR2_X1 i_0_263 (.ZN (n_0_141), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_262 (.ZN (u[60]), .A (y[60]), .B (n_0_141));
XNOR2_X1 i_0_261 (.ZN (n_0_140), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_260 (.ZN (u[59]), .A (y[59]), .B (n_0_140));
XNOR2_X1 i_0_259 (.ZN (n_0_139), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_258 (.ZN (u[58]), .A (y[58]), .B (n_0_139));
XNOR2_X1 i_0_257 (.ZN (n_0_138), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_256 (.ZN (u[57]), .A (y[57]), .B (n_0_138));
XNOR2_X1 i_0_255 (.ZN (n_0_137), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_254 (.ZN (u[56]), .A (y[56]), .B (n_0_137));
XNOR2_X1 i_0_253 (.ZN (n_0_136), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_252 (.ZN (u[55]), .A (y[55]), .B (n_0_136));
XNOR2_X1 i_0_251 (.ZN (n_0_135), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_250 (.ZN (u[54]), .A (y[54]), .B (n_0_135));
XNOR2_X1 i_0_249 (.ZN (n_0_134), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_248 (.ZN (u[53]), .A (y[53]), .B (n_0_134));
XNOR2_X1 i_0_247 (.ZN (n_0_133), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_246 (.ZN (u[52]), .A (y[52]), .B (n_0_133));
XNOR2_X1 i_0_245 (.ZN (n_0_132), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_244 (.ZN (u[51]), .A (y[51]), .B (n_0_132));
XNOR2_X1 i_0_243 (.ZN (n_0_131), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_242 (.ZN (u[50]), .A (y[50]), .B (n_0_131));
XNOR2_X1 i_0_241 (.ZN (n_0_130), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_240 (.ZN (u[49]), .A (y[49]), .B (n_0_130));
XNOR2_X1 i_0_239 (.ZN (n_0_129), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_238 (.ZN (u[48]), .A (y[48]), .B (n_0_129));
XNOR2_X1 i_0_237 (.ZN (n_0_128), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_236 (.ZN (u[47]), .A (y[47]), .B (n_0_128));
XNOR2_X1 i_0_235 (.ZN (n_0_127), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_234 (.ZN (u[46]), .A (y[46]), .B (n_0_127));
XNOR2_X1 i_0_233 (.ZN (n_0_126), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_232 (.ZN (u[45]), .A (y[45]), .B (n_0_126));
XNOR2_X1 i_0_231 (.ZN (n_0_125), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_230 (.ZN (u[44]), .A (y[44]), .B (n_0_125));
XNOR2_X1 i_0_229 (.ZN (n_0_124), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_228 (.ZN (u[43]), .A (y[43]), .B (n_0_124));
XNOR2_X1 i_0_227 (.ZN (n_0_123), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_226 (.ZN (u[42]), .A (y[42]), .B (n_0_123));
XNOR2_X1 i_0_225 (.ZN (n_0_122), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_224 (.ZN (u[41]), .A (y[41]), .B (n_0_122));
XNOR2_X1 i_0_223 (.ZN (n_0_121), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_222 (.ZN (u[40]), .A (y[40]), .B (n_0_121));
XNOR2_X1 i_0_221 (.ZN (n_0_120), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_220 (.ZN (u[39]), .A (y[39]), .B (n_0_120));
XNOR2_X1 i_0_219 (.ZN (n_0_119), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_218 (.ZN (u[38]), .A (y[38]), .B (n_0_119));
XNOR2_X1 i_0_217 (.ZN (n_0_118), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_216 (.ZN (u[37]), .A (y[37]), .B (n_0_118));
XNOR2_X1 i_0_215 (.ZN (n_0_117), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_214 (.ZN (u[36]), .A (y[36]), .B (n_0_117));
XNOR2_X1 i_0_213 (.ZN (n_0_116), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_212 (.ZN (u[35]), .A (y[35]), .B (n_0_116));
XNOR2_X1 i_0_211 (.ZN (n_0_115), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_210 (.ZN (u[34]), .A (y[34]), .B (n_0_115));
XNOR2_X1 i_0_209 (.ZN (n_0_114), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_208 (.ZN (u[33]), .A (y[33]), .B (n_0_114));
XNOR2_X1 i_0_207 (.ZN (n_0_113), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_206 (.ZN (u[32]), .A (y[32]), .B (n_0_113));
XNOR2_X1 i_0_205 (.ZN (n_0_112), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_204 (.ZN (u[31]), .A (y[31]), .B (n_0_112));
XNOR2_X1 i_0_203 (.ZN (n_0_111), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_202 (.ZN (u[30]), .A (y[30]), .B (n_0_111));
XNOR2_X1 i_0_201 (.ZN (n_0_110), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_200 (.ZN (u[29]), .A (y[29]), .B (n_0_110));
XNOR2_X1 i_0_199 (.ZN (n_0_109), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_198 (.ZN (u[28]), .A (y[28]), .B (n_0_109));
XNOR2_X1 i_0_197 (.ZN (n_0_108), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_196 (.ZN (u[27]), .A (y[27]), .B (n_0_108));
XNOR2_X1 i_0_195 (.ZN (n_0_107), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_194 (.ZN (u[26]), .A (y[26]), .B (n_0_107));
XNOR2_X1 i_0_193 (.ZN (n_0_106), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_192 (.ZN (u[25]), .A (y[25]), .B (n_0_106));
XNOR2_X1 i_0_191 (.ZN (n_0_105), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_190 (.ZN (u[24]), .A (y[24]), .B (n_0_105));
XNOR2_X1 i_0_189 (.ZN (n_0_104), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_188 (.ZN (u[23]), .A (y[23]), .B (n_0_104));
XNOR2_X1 i_0_187 (.ZN (n_0_103), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_186 (.ZN (u[22]), .A (y[22]), .B (n_0_103));
XNOR2_X1 i_0_185 (.ZN (n_0_102), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_184 (.ZN (u[21]), .A (y[21]), .B (n_0_102));
XNOR2_X1 i_0_183 (.ZN (n_0_101), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_182 (.ZN (u[20]), .A (y[20]), .B (n_0_101));
XNOR2_X1 i_0_181 (.ZN (n_0_100), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_180 (.ZN (u[19]), .A (y[19]), .B (n_0_100));
XNOR2_X1 i_0_179 (.ZN (n_0_99), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_178 (.ZN (u[18]), .A (y[18]), .B (n_0_99));
XNOR2_X1 i_0_177 (.ZN (n_0_98), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_176 (.ZN (u[17]), .A (y[17]), .B (n_0_98));
XNOR2_X1 i_0_175 (.ZN (n_0_97), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_174 (.ZN (u[16]), .A (y[16]), .B (n_0_97));
XNOR2_X2 i_0_173 (.ZN (n_0_96), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_172 (.ZN (u[15]), .A (y[15]), .B (n_0_96));
XOR2_X2 i_0_171 (.Z (u[14]), .A (y[14]), .B (x[14]));
XOR2_X2 i_0_170 (.Z (u[13]), .A (y[13]), .B (x[13]));
XOR2_X2 i_0_169 (.Z (u[12]), .A (y[12]), .B (x[12]));
XOR2_X2 i_0_166 (.Z (u[9]), .A (x[9]), .B (y[9]));
XOR2_X2 i_0_165 (.Z (u[8]), .A (y[8]), .B (x[8]));
XOR2_X2 i_0_164 (.Z (u[7]), .A (y[7]), .B (x[7]));
XOR2_X1 i_0_163 (.Z (u[6]), .A (y[6]), .B (x[6]));
NAND2_X1 i_0_157 (.ZN (n_0_95), .A1 (z[62]), .A2 (x[62]));
OAI21_X1 i_0_156 (.ZN (n_0_94), .A (y[62]), .B1 (z[62]), .B2 (x[62]));
NAND2_X1 i_0_155 (.ZN (v[63]), .A1 (n_0_95), .A2 (n_0_94));
NAND2_X1 i_0_154 (.ZN (n_0_93), .A1 (z[61]), .A2 (x[61]));
OAI21_X1 i_0_153 (.ZN (n_0_92), .A (y[61]), .B1 (z[61]), .B2 (x[61]));
NAND2_X1 i_0_152 (.ZN (v[62]), .A1 (n_0_93), .A2 (n_0_92));
NAND2_X1 i_0_151 (.ZN (n_0_91), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_150 (.ZN (n_0_90), .A (y[60]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_149 (.ZN (v[61]), .A1 (n_0_91), .A2 (n_0_90));
NAND2_X1 i_0_148 (.ZN (n_0_89), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_147 (.ZN (n_0_88), .A (y[59]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_146 (.ZN (v[60]), .A1 (n_0_89), .A2 (n_0_88));
NAND2_X1 i_0_145 (.ZN (n_0_87), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_144 (.ZN (n_0_86), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_143 (.ZN (v[59]), .A1 (n_0_87), .A2 (n_0_86));
NAND2_X1 i_0_142 (.ZN (n_0_85), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_141 (.ZN (n_0_84), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_140 (.ZN (v[58]), .A1 (n_0_85), .A2 (n_0_84));
NAND2_X1 i_0_139 (.ZN (n_0_83), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_138 (.ZN (n_0_82), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_137 (.ZN (v[57]), .A1 (n_0_83), .A2 (n_0_82));
NAND2_X1 i_0_136 (.ZN (n_0_81), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_135 (.ZN (n_0_80), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_134 (.ZN (v[56]), .A1 (n_0_81), .A2 (n_0_80));
NAND2_X1 i_0_133 (.ZN (n_0_79), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_132 (.ZN (n_0_78), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_131 (.ZN (v[55]), .A1 (n_0_79), .A2 (n_0_78));
NAND2_X1 i_0_130 (.ZN (n_0_77), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_129 (.ZN (n_0_76), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_128 (.ZN (v[54]), .A1 (n_0_77), .A2 (n_0_76));
NAND2_X1 i_0_127 (.ZN (n_0_75), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_126 (.ZN (n_0_74), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_125 (.ZN (v[53]), .A1 (n_0_75), .A2 (n_0_74));
NAND2_X1 i_0_124 (.ZN (n_0_73), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_123 (.ZN (n_0_72), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_122 (.ZN (v[52]), .A1 (n_0_73), .A2 (n_0_72));
NAND2_X1 i_0_121 (.ZN (n_0_71), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_120 (.ZN (n_0_70), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_119 (.ZN (v[51]), .A1 (n_0_71), .A2 (n_0_70));
NAND2_X1 i_0_118 (.ZN (n_0_69), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_117 (.ZN (n_0_68), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_116 (.ZN (v[50]), .A1 (n_0_69), .A2 (n_0_68));
NAND2_X1 i_0_115 (.ZN (n_0_67), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_114 (.ZN (n_0_66), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_113 (.ZN (v[49]), .A1 (n_0_67), .A2 (n_0_66));
NAND2_X1 i_0_112 (.ZN (n_0_65), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_111 (.ZN (n_0_64), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_110 (.ZN (v[48]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_109 (.ZN (n_0_63), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_108 (.ZN (n_0_62), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_107 (.ZN (v[47]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_106 (.ZN (n_0_61), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_105 (.ZN (n_0_60), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_104 (.ZN (v[46]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_103 (.ZN (n_0_59), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_102 (.ZN (n_0_58), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_101 (.ZN (v[45]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_100 (.ZN (n_0_57), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_99 (.ZN (n_0_56), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_98 (.ZN (v[44]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_97 (.ZN (n_0_55), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_96 (.ZN (n_0_54), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_95 (.ZN (v[43]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_94 (.ZN (n_0_53), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_93 (.ZN (n_0_52), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_92 (.ZN (v[42]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_91 (.ZN (n_0_51), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_90 (.ZN (n_0_50), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_89 (.ZN (v[41]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_88 (.ZN (n_0_49), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_87 (.ZN (n_0_48), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_86 (.ZN (v[40]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_85 (.ZN (n_0_47), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_84 (.ZN (n_0_46), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_83 (.ZN (v[39]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_82 (.ZN (n_0_45), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_81 (.ZN (n_0_44), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_80 (.ZN (v[38]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_79 (.ZN (n_0_43), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_78 (.ZN (n_0_42), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_77 (.ZN (v[37]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_76 (.ZN (n_0_41), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_75 (.ZN (n_0_40), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_74 (.ZN (v[36]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_73 (.ZN (n_0_39), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_72 (.ZN (n_0_38), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_71 (.ZN (v[35]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_70 (.ZN (n_0_37), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_69 (.ZN (n_0_36), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_68 (.ZN (v[34]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_67 (.ZN (n_0_35), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_66 (.ZN (n_0_34), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_65 (.ZN (v[33]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_64 (.ZN (n_0_33), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_63 (.ZN (n_0_32), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_62 (.ZN (v[32]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_61 (.ZN (n_0_31), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_60 (.ZN (n_0_30), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_59 (.ZN (v[31]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_58 (.ZN (n_0_29), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_57 (.ZN (n_0_28), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_56 (.ZN (v[30]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_55 (.ZN (n_0_27), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_54 (.ZN (n_0_26), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_53 (.ZN (v[29]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_52 (.ZN (n_0_25), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_51 (.ZN (n_0_24), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_50 (.ZN (v[28]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_49 (.ZN (n_0_23), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_48 (.ZN (n_0_22), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_47 (.ZN (v[27]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_46 (.ZN (n_0_21), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_45 (.ZN (n_0_20), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_44 (.ZN (v[26]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_43 (.ZN (n_0_19), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_42 (.ZN (n_0_18), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_41 (.ZN (v[25]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_40 (.ZN (n_0_17), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_39 (.ZN (n_0_16), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_38 (.ZN (v[24]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_37 (.ZN (n_0_15), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_36 (.ZN (n_0_14), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_35 (.ZN (v[23]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_34 (.ZN (n_0_13), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_33 (.ZN (n_0_12), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_32 (.ZN (v[22]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_31 (.ZN (n_0_11), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_30 (.ZN (n_0_10), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_29 (.ZN (v[21]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_28 (.ZN (n_0_9), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_27 (.ZN (n_0_8), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_26 (.ZN (v[20]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_25 (.ZN (n_0_7), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_24 (.ZN (n_0_6), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_23 (.ZN (v[19]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_22 (.ZN (n_0_5), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_21 (.ZN (n_0_4), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_20 (.ZN (v[18]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_19 (.ZN (n_0_3), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_18 (.ZN (n_0_2), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_17 (.ZN (v[17]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_16 (.ZN (n_0_1), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_15 (.ZN (n_0_0), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_14 (.ZN (v[16]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_13 (.ZN (v[15]), .A1 (y[14]), .A2 (x[14]));
AND2_X1 i_0_12 (.ZN (v[14]), .A1 (y[13]), .A2 (x[13]));
AND2_X2 i_0_11 (.ZN (v[13]), .A1 (y[12]), .A2 (x[12]));
AND2_X1 i_0_10 (.ZN (v[12]), .A1 (y[11]), .A2 (x[11]));
AND2_X1 i_0_9 (.ZN (v[11]), .A1 (y[10]), .A2 (x[10]));
AND2_X2 i_0_8 (.ZN (v[10]), .A1 (y[9]), .A2 (x[9]));
AND2_X2 i_0_7 (.ZN (v[9]), .A1 (y[8]), .A2 (x[8]));
AND2_X2 i_0_6 (.ZN (v[8]), .A1 (y[7]), .A2 (x[7]));
AND2_X2 i_0_5 (.ZN (v[7]), .A1 (y[6]), .A2 (x[6]));
INV_X1 slo__mro_c8 (.ZN (slo__mro_n9), .A (y[11]));
XNOR2_X2 slo__mro_c9 (.ZN (u[11]), .A (x[11]), .B (slo__mro_n9));

endmodule //CSA__5_206

module CSA__5_203 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;


XNOR2_X1 i_0_199 (.ZN (n_0_114), .A (z[63]), .B (x[63]));
XNOR2_X1 i_0_198 (.ZN (u[63]), .A (y[63]), .B (n_0_114));
XNOR2_X1 i_0_197 (.ZN (n_0_113), .A (z[62]), .B (x[62]));
XNOR2_X1 i_0_196 (.ZN (u[62]), .A (y[62]), .B (n_0_113));
XNOR2_X1 i_0_195 (.ZN (n_0_112), .A (z[61]), .B (x[61]));
XNOR2_X1 i_0_194 (.ZN (u[61]), .A (y[61]), .B (n_0_112));
XNOR2_X1 i_0_193 (.ZN (n_0_111), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_192 (.ZN (u[60]), .A (y[60]), .B (n_0_111));
XNOR2_X1 i_0_191 (.ZN (n_0_110), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_190 (.ZN (u[59]), .A (y[59]), .B (n_0_110));
XNOR2_X1 i_0_189 (.ZN (n_0_109), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_188 (.ZN (u[58]), .A (y[58]), .B (n_0_109));
XNOR2_X1 i_0_187 (.ZN (n_0_108), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_186 (.ZN (u[57]), .A (y[57]), .B (n_0_108));
XNOR2_X1 i_0_185 (.ZN (n_0_107), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_184 (.ZN (u[56]), .A (y[56]), .B (n_0_107));
XNOR2_X1 i_0_183 (.ZN (n_0_106), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_182 (.ZN (u[55]), .A (y[55]), .B (n_0_106));
XNOR2_X1 i_0_181 (.ZN (n_0_105), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_180 (.ZN (u[54]), .A (y[54]), .B (n_0_105));
XNOR2_X1 i_0_179 (.ZN (n_0_104), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_178 (.ZN (u[53]), .A (y[53]), .B (n_0_104));
XNOR2_X1 i_0_177 (.ZN (n_0_103), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_176 (.ZN (u[52]), .A (y[52]), .B (n_0_103));
XNOR2_X1 i_0_175 (.ZN (n_0_102), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_174 (.ZN (u[51]), .A (y[51]), .B (n_0_102));
XNOR2_X1 i_0_173 (.ZN (n_0_101), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_172 (.ZN (u[50]), .A (y[50]), .B (n_0_101));
XNOR2_X1 i_0_171 (.ZN (n_0_100), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_170 (.ZN (u[49]), .A (y[49]), .B (n_0_100));
XNOR2_X1 i_0_169 (.ZN (n_0_99), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_168 (.ZN (u[48]), .A (y[48]), .B (n_0_99));
XNOR2_X1 i_0_167 (.ZN (n_0_98), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_166 (.ZN (u[47]), .A (y[47]), .B (n_0_98));
XNOR2_X1 i_0_165 (.ZN (n_0_97), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_164 (.ZN (u[46]), .A (y[46]), .B (n_0_97));
XNOR2_X1 i_0_163 (.ZN (n_0_96), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_162 (.ZN (u[45]), .A (y[45]), .B (n_0_96));
XNOR2_X1 i_0_161 (.ZN (n_0_95), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_160 (.ZN (u[44]), .A (y[44]), .B (n_0_95));
XNOR2_X1 i_0_159 (.ZN (n_0_94), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_158 (.ZN (u[43]), .A (y[43]), .B (n_0_94));
XNOR2_X1 i_0_157 (.ZN (n_0_93), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_156 (.ZN (u[42]), .A (y[42]), .B (n_0_93));
XNOR2_X1 i_0_155 (.ZN (n_0_92), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_154 (.ZN (u[41]), .A (y[41]), .B (n_0_92));
XNOR2_X1 i_0_153 (.ZN (n_0_91), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_152 (.ZN (u[40]), .A (y[40]), .B (n_0_91));
XNOR2_X1 i_0_151 (.ZN (n_0_90), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_150 (.ZN (u[39]), .A (y[39]), .B (n_0_90));
XNOR2_X1 i_0_149 (.ZN (n_0_89), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_148 (.ZN (u[38]), .A (y[38]), .B (n_0_89));
XNOR2_X1 i_0_147 (.ZN (n_0_88), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_146 (.ZN (u[37]), .A (y[37]), .B (n_0_88));
XNOR2_X1 i_0_145 (.ZN (n_0_87), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_144 (.ZN (u[36]), .A (y[36]), .B (n_0_87));
XNOR2_X1 i_0_143 (.ZN (n_0_86), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_142 (.ZN (u[35]), .A (y[35]), .B (n_0_86));
XNOR2_X1 i_0_141 (.ZN (n_0_85), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_140 (.ZN (u[34]), .A (y[34]), .B (n_0_85));
XNOR2_X1 i_0_139 (.ZN (n_0_84), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_138 (.ZN (u[33]), .A (y[33]), .B (n_0_84));
XNOR2_X1 i_0_137 (.ZN (n_0_83), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_136 (.ZN (u[32]), .A (y[32]), .B (n_0_83));
XNOR2_X1 i_0_135 (.ZN (n_0_82), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_134 (.ZN (u[31]), .A (y[31]), .B (n_0_82));
XNOR2_X1 i_0_133 (.ZN (n_0_81), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_132 (.ZN (u[30]), .A (y[30]), .B (n_0_81));
XNOR2_X1 i_0_131 (.ZN (n_0_80), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_130 (.ZN (u[29]), .A (y[29]), .B (n_0_80));
XNOR2_X1 i_0_129 (.ZN (n_0_79), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_128 (.ZN (u[28]), .A (y[28]), .B (n_0_79));
XNOR2_X1 i_0_127 (.ZN (n_0_78), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_126 (.ZN (u[27]), .A (y[27]), .B (n_0_78));
XNOR2_X1 i_0_125 (.ZN (n_0_77), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_124 (.ZN (u[26]), .A (y[26]), .B (n_0_77));
XNOR2_X1 i_0_123 (.ZN (n_0_76), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_122 (.ZN (u[25]), .A (y[25]), .B (n_0_76));
XOR2_X1 i_0_121 (.Z (u[24]), .A (y[24]), .B (x[24]));
XOR2_X1 i_0_120 (.Z (u[23]), .A (y[23]), .B (x[23]));
XOR2_X1 i_0_119 (.Z (u[22]), .A (y[22]), .B (x[22]));
XOR2_X1 i_0_118 (.Z (u[21]), .A (y[21]), .B (x[21]));
NAND2_X1 i_0_117 (.ZN (n_0_75), .A1 (z[62]), .A2 (x[62]));
OAI21_X1 i_0_116 (.ZN (n_0_74), .A (y[62]), .B1 (z[62]), .B2 (x[62]));
NAND2_X1 i_0_115 (.ZN (v[63]), .A1 (n_0_75), .A2 (n_0_74));
NAND2_X1 i_0_114 (.ZN (n_0_73), .A1 (z[61]), .A2 (x[61]));
OAI21_X1 i_0_113 (.ZN (n_0_72), .A (y[61]), .B1 (z[61]), .B2 (x[61]));
NAND2_X1 i_0_112 (.ZN (v[62]), .A1 (n_0_73), .A2 (n_0_72));
NAND2_X1 i_0_111 (.ZN (n_0_71), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_110 (.ZN (n_0_70), .A (y[60]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_109 (.ZN (v[61]), .A1 (n_0_71), .A2 (n_0_70));
NAND2_X1 i_0_108 (.ZN (n_0_69), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_107 (.ZN (n_0_68), .A (y[59]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_106 (.ZN (v[60]), .A1 (n_0_69), .A2 (n_0_68));
NAND2_X1 i_0_105 (.ZN (n_0_67), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_104 (.ZN (n_0_66), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_103 (.ZN (v[59]), .A1 (n_0_67), .A2 (n_0_66));
NAND2_X1 i_0_102 (.ZN (n_0_65), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_101 (.ZN (n_0_64), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_100 (.ZN (v[58]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_99 (.ZN (n_0_63), .A1 (y[56]), .A2 (z[56]));
OAI21_X1 i_0_98 (.ZN (n_0_62), .A (x[56]), .B1 (z[56]), .B2 (y[56]));
NAND2_X1 i_0_97 (.ZN (v[57]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_96 (.ZN (n_0_61), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_95 (.ZN (n_0_60), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_94 (.ZN (v[56]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_93 (.ZN (n_0_59), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_92 (.ZN (n_0_58), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_91 (.ZN (v[55]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_90 (.ZN (n_0_57), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_89 (.ZN (n_0_56), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_88 (.ZN (v[54]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_87 (.ZN (n_0_55), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_86 (.ZN (n_0_54), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_85 (.ZN (v[53]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_84 (.ZN (n_0_53), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_83 (.ZN (n_0_52), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_82 (.ZN (v[52]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_81 (.ZN (n_0_51), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_80 (.ZN (n_0_50), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_79 (.ZN (v[51]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_78 (.ZN (n_0_49), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_77 (.ZN (n_0_48), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_76 (.ZN (v[50]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_75 (.ZN (n_0_47), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_74 (.ZN (n_0_46), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_73 (.ZN (v[49]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_72 (.ZN (n_0_45), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_71 (.ZN (n_0_44), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_70 (.ZN (v[48]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_69 (.ZN (n_0_43), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_68 (.ZN (n_0_42), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_67 (.ZN (v[47]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_66 (.ZN (n_0_41), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_65 (.ZN (n_0_40), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_64 (.ZN (v[46]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_63 (.ZN (n_0_39), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_62 (.ZN (n_0_38), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_61 (.ZN (v[45]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_60 (.ZN (n_0_37), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_59 (.ZN (n_0_36), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_58 (.ZN (v[44]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_57 (.ZN (n_0_35), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_56 (.ZN (n_0_34), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_55 (.ZN (v[43]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_54 (.ZN (n_0_33), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_53 (.ZN (n_0_32), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_52 (.ZN (v[42]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_51 (.ZN (n_0_31), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_50 (.ZN (n_0_30), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_49 (.ZN (v[41]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_48 (.ZN (n_0_29), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_47 (.ZN (n_0_28), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_46 (.ZN (v[40]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_45 (.ZN (n_0_27), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_44 (.ZN (n_0_26), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_43 (.ZN (v[39]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_42 (.ZN (n_0_25), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_41 (.ZN (n_0_24), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_40 (.ZN (v[38]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_39 (.ZN (n_0_23), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_38 (.ZN (n_0_22), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_37 (.ZN (v[37]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_36 (.ZN (n_0_21), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_35 (.ZN (n_0_20), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_34 (.ZN (v[36]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_33 (.ZN (n_0_19), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_32 (.ZN (n_0_18), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_31 (.ZN (v[35]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_30 (.ZN (n_0_17), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_29 (.ZN (n_0_16), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_28 (.ZN (v[34]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_27 (.ZN (n_0_15), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_26 (.ZN (n_0_14), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_25 (.ZN (v[33]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_24 (.ZN (n_0_13), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_23 (.ZN (n_0_12), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_22 (.ZN (v[32]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_21 (.ZN (n_0_11), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_20 (.ZN (n_0_10), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_19 (.ZN (v[31]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_18 (.ZN (n_0_9), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_17 (.ZN (n_0_8), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_16 (.ZN (v[30]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_15 (.ZN (n_0_7), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_14 (.ZN (n_0_6), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_13 (.ZN (v[29]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_12 (.ZN (n_0_5), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_11 (.ZN (n_0_4), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_10 (.ZN (v[28]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_9 (.ZN (n_0_3), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_8 (.ZN (n_0_2), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_7 (.ZN (v[27]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_6 (.ZN (n_0_1), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_5 (.ZN (n_0_0), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_4 (.ZN (v[26]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_3 (.ZN (v[25]), .A1 (y[24]), .A2 (x[24]));
AND2_X1 i_0_2 (.ZN (v[24]), .A1 (y[23]), .A2 (x[23]));
AND2_X1 i_0_1 (.ZN (v[23]), .A1 (y[22]), .A2 (x[22]));
AND2_X1 i_0_0 (.ZN (v[22]), .A1 (y[21]), .A2 (x[21]));

endmodule //CSA__5_203

module CSA__5_200 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;


XNOR2_X1 i_0_231 (.ZN (n_0_108), .A (z[63]), .B (x[63]));
XNOR2_X1 i_0_230 (.ZN (u[63]), .A (y[63]), .B (n_0_108));
XNOR2_X1 i_0_229 (.ZN (n_0_107), .A (z[62]), .B (x[62]));
XNOR2_X1 i_0_228 (.ZN (u[62]), .A (y[63]), .B (n_0_107));
XNOR2_X1 i_0_227 (.ZN (n_0_106), .A (z[61]), .B (x[61]));
XNOR2_X1 i_0_226 (.ZN (u[61]), .A (y[63]), .B (n_0_106));
XNOR2_X1 i_0_225 (.ZN (n_0_105), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_224 (.ZN (u[60]), .A (y[63]), .B (n_0_105));
XNOR2_X1 i_0_223 (.ZN (n_0_104), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_222 (.ZN (u[59]), .A (y[59]), .B (n_0_104));
XNOR2_X1 i_0_221 (.ZN (n_0_103), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_220 (.ZN (u[58]), .A (y[58]), .B (n_0_103));
XNOR2_X1 i_0_219 (.ZN (n_0_102), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_218 (.ZN (u[57]), .A (y[57]), .B (n_0_102));
XNOR2_X1 i_0_217 (.ZN (n_0_101), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_216 (.ZN (u[56]), .A (y[56]), .B (n_0_101));
XNOR2_X1 i_0_215 (.ZN (n_0_100), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_214 (.ZN (u[55]), .A (y[55]), .B (n_0_100));
XNOR2_X1 i_0_213 (.ZN (n_0_99), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_212 (.ZN (u[54]), .A (y[54]), .B (n_0_99));
XNOR2_X1 i_0_211 (.ZN (n_0_98), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_210 (.ZN (u[53]), .A (y[53]), .B (n_0_98));
XNOR2_X1 i_0_209 (.ZN (n_0_97), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_208 (.ZN (u[52]), .A (y[52]), .B (n_0_97));
XNOR2_X1 i_0_207 (.ZN (n_0_96), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_206 (.ZN (u[51]), .A (y[51]), .B (n_0_96));
XNOR2_X1 i_0_205 (.ZN (n_0_95), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_204 (.ZN (u[50]), .A (y[50]), .B (n_0_95));
XNOR2_X1 i_0_203 (.ZN (n_0_94), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_202 (.ZN (u[49]), .A (y[49]), .B (n_0_94));
XNOR2_X1 i_0_201 (.ZN (n_0_93), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_200 (.ZN (u[48]), .A (y[48]), .B (n_0_93));
XNOR2_X1 i_0_199 (.ZN (n_0_92), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_198 (.ZN (u[47]), .A (y[47]), .B (n_0_92));
XNOR2_X1 i_0_197 (.ZN (n_0_91), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_196 (.ZN (u[46]), .A (y[46]), .B (n_0_91));
XNOR2_X1 i_0_195 (.ZN (n_0_90), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_194 (.ZN (u[45]), .A (y[45]), .B (n_0_90));
XNOR2_X1 i_0_193 (.ZN (n_0_89), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_192 (.ZN (u[44]), .A (y[44]), .B (n_0_89));
XNOR2_X1 i_0_191 (.ZN (n_0_88), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_190 (.ZN (u[43]), .A (y[43]), .B (n_0_88));
XNOR2_X1 i_0_189 (.ZN (n_0_87), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_188 (.ZN (u[42]), .A (y[42]), .B (n_0_87));
XNOR2_X1 i_0_187 (.ZN (n_0_86), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_186 (.ZN (u[41]), .A (y[41]), .B (n_0_86));
XNOR2_X1 i_0_185 (.ZN (n_0_85), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_184 (.ZN (u[40]), .A (y[40]), .B (n_0_85));
XNOR2_X1 i_0_183 (.ZN (n_0_84), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_182 (.ZN (u[39]), .A (y[39]), .B (n_0_84));
XNOR2_X1 i_0_181 (.ZN (n_0_83), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_180 (.ZN (u[38]), .A (y[38]), .B (n_0_83));
XNOR2_X1 i_0_179 (.ZN (n_0_82), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_178 (.ZN (u[37]), .A (y[37]), .B (n_0_82));
XNOR2_X1 i_0_177 (.ZN (n_0_81), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_176 (.ZN (u[36]), .A (y[36]), .B (n_0_81));
XNOR2_X1 i_0_175 (.ZN (n_0_80), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_174 (.ZN (u[35]), .A (y[35]), .B (n_0_80));
XNOR2_X1 i_0_173 (.ZN (n_0_79), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_172 (.ZN (u[34]), .A (y[34]), .B (n_0_79));
XNOR2_X1 i_0_171 (.ZN (n_0_78), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_170 (.ZN (u[33]), .A (y[33]), .B (n_0_78));
XNOR2_X1 i_0_169 (.ZN (n_0_77), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_168 (.ZN (u[32]), .A (y[32]), .B (n_0_77));
XNOR2_X1 i_0_167 (.ZN (n_0_76), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_166 (.ZN (u[31]), .A (y[31]), .B (n_0_76));
XNOR2_X1 i_0_165 (.ZN (n_0_75), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_164 (.ZN (u[30]), .A (y[30]), .B (n_0_75));
XNOR2_X1 i_0_163 (.ZN (n_0_74), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_162 (.ZN (u[29]), .A (y[29]), .B (n_0_74));
XNOR2_X1 i_0_161 (.ZN (n_0_73), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_160 (.ZN (u[28]), .A (y[28]), .B (n_0_73));
XNOR2_X1 i_0_159 (.ZN (n_0_72), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_158 (.ZN (u[27]), .A (y[27]), .B (n_0_72));
XOR2_X1 i_0_157 (.Z (u[26]), .A (y[26]), .B (x[26]));
XOR2_X1 i_0_156 (.Z (u[25]), .A (y[25]), .B (x[25]));
XOR2_X1 i_0_155 (.Z (u[24]), .A (y[24]), .B (x[24]));
NAND2_X1 i_0_132 (.ZN (n_0_71), .A1 (z[62]), .A2 (x[62]));
OAI21_X1 i_0_131 (.ZN (n_0_70), .A (y[63]), .B1 (z[62]), .B2 (x[62]));
NAND2_X1 i_0_130 (.ZN (v[63]), .A1 (n_0_71), .A2 (n_0_70));
NAND2_X1 i_0_129 (.ZN (n_0_69), .A1 (z[61]), .A2 (x[61]));
OAI21_X1 i_0_128 (.ZN (n_0_68), .A (y[63]), .B1 (z[61]), .B2 (x[61]));
NAND2_X1 i_0_127 (.ZN (v[62]), .A1 (n_0_69), .A2 (n_0_68));
NAND2_X1 i_0_126 (.ZN (n_0_67), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_125 (.ZN (n_0_66), .A (y[63]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_124 (.ZN (v[61]), .A1 (n_0_67), .A2 (n_0_66));
NAND2_X1 i_0_123 (.ZN (n_0_65), .A1 (y[59]), .A2 (z[59]));
OAI21_X1 i_0_122 (.ZN (n_0_64), .A (x[59]), .B1 (z[59]), .B2 (y[59]));
NAND2_X1 i_0_121 (.ZN (v[60]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_120 (.ZN (n_0_63), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_119 (.ZN (n_0_62), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_118 (.ZN (v[59]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_117 (.ZN (n_0_61), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_116 (.ZN (n_0_60), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_115 (.ZN (v[58]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_114 (.ZN (n_0_59), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_113 (.ZN (n_0_58), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_112 (.ZN (v[57]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_111 (.ZN (n_0_57), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_110 (.ZN (n_0_56), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_109 (.ZN (v[56]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_108 (.ZN (n_0_55), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_107 (.ZN (n_0_54), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_106 (.ZN (v[55]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_105 (.ZN (n_0_53), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_104 (.ZN (n_0_52), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_103 (.ZN (v[54]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_102 (.ZN (n_0_51), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_101 (.ZN (n_0_50), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_100 (.ZN (v[53]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_99 (.ZN (n_0_49), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_98 (.ZN (n_0_48), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_97 (.ZN (v[52]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_96 (.ZN (n_0_47), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_95 (.ZN (n_0_46), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_94 (.ZN (v[51]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_93 (.ZN (n_0_45), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_92 (.ZN (n_0_44), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_91 (.ZN (v[50]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_90 (.ZN (n_0_43), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_89 (.ZN (n_0_42), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_88 (.ZN (v[49]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_87 (.ZN (n_0_41), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_86 (.ZN (n_0_40), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_85 (.ZN (v[48]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_84 (.ZN (n_0_39), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_83 (.ZN (n_0_38), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_82 (.ZN (v[47]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_81 (.ZN (n_0_37), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_80 (.ZN (n_0_36), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_79 (.ZN (v[46]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_78 (.ZN (n_0_35), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_77 (.ZN (n_0_34), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_76 (.ZN (v[45]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_75 (.ZN (n_0_33), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_74 (.ZN (n_0_32), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_73 (.ZN (v[44]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_72 (.ZN (n_0_31), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_71 (.ZN (n_0_30), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_70 (.ZN (v[43]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_69 (.ZN (n_0_29), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_68 (.ZN (n_0_28), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_67 (.ZN (v[42]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_66 (.ZN (n_0_27), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_65 (.ZN (n_0_26), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_64 (.ZN (v[41]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_63 (.ZN (n_0_25), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_62 (.ZN (n_0_24), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_61 (.ZN (v[40]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_60 (.ZN (n_0_23), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_59 (.ZN (n_0_22), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_58 (.ZN (v[39]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_57 (.ZN (n_0_21), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_56 (.ZN (n_0_20), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_55 (.ZN (v[38]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_54 (.ZN (n_0_19), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_53 (.ZN (n_0_18), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_52 (.ZN (v[37]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_51 (.ZN (n_0_17), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_50 (.ZN (n_0_16), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_49 (.ZN (v[36]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_48 (.ZN (n_0_15), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_47 (.ZN (n_0_14), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_46 (.ZN (v[35]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_45 (.ZN (n_0_13), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_44 (.ZN (n_0_12), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_43 (.ZN (v[34]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_42 (.ZN (n_0_11), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_41 (.ZN (n_0_10), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_40 (.ZN (v[33]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_39 (.ZN (n_0_9), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_38 (.ZN (n_0_8), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_37 (.ZN (v[32]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_36 (.ZN (n_0_7), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_35 (.ZN (n_0_6), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_34 (.ZN (v[31]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_33 (.ZN (n_0_5), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_32 (.ZN (n_0_4), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_31 (.ZN (v[30]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_30 (.ZN (n_0_3), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_29 (.ZN (n_0_2), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_28 (.ZN (v[29]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_27 (.ZN (n_0_1), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_26 (.ZN (n_0_0), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_25 (.ZN (v[28]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_24 (.ZN (v[27]), .A1 (y[26]), .A2 (x[26]));
AND2_X1 i_0_23 (.ZN (v[26]), .A1 (y[25]), .A2 (x[25]));
AND2_X1 i_0_22 (.ZN (v[25]), .A1 (y[24]), .A2 (x[24]));

endmodule //CSA__5_200

module CSA__5_197 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;


XNOR2_X1 i_0_163 (.ZN (n_0_96), .A (z[63]), .B (x[63]));
XNOR2_X1 i_0_162 (.ZN (u[63]), .A (y[63]), .B (n_0_96));
XNOR2_X1 i_0_161 (.ZN (n_0_95), .A (z[63]), .B (x[62]));
XNOR2_X1 i_0_160 (.ZN (u[62]), .A (y[62]), .B (n_0_95));
XNOR2_X1 i_0_159 (.ZN (n_0_94), .A (z[61]), .B (x[61]));
XNOR2_X1 i_0_158 (.ZN (u[61]), .A (y[61]), .B (n_0_94));
XNOR2_X1 i_0_157 (.ZN (n_0_93), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_156 (.ZN (u[60]), .A (y[60]), .B (n_0_93));
XNOR2_X1 i_0_155 (.ZN (n_0_92), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_154 (.ZN (u[59]), .A (y[59]), .B (n_0_92));
XNOR2_X1 i_0_153 (.ZN (n_0_91), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_152 (.ZN (u[58]), .A (y[58]), .B (n_0_91));
XNOR2_X1 i_0_151 (.ZN (n_0_90), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_150 (.ZN (u[57]), .A (y[57]), .B (n_0_90));
XNOR2_X1 i_0_149 (.ZN (n_0_89), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_148 (.ZN (u[56]), .A (y[56]), .B (n_0_89));
XNOR2_X1 i_0_147 (.ZN (n_0_88), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_146 (.ZN (u[55]), .A (y[55]), .B (n_0_88));
XNOR2_X1 i_0_145 (.ZN (n_0_87), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_144 (.ZN (u[54]), .A (y[54]), .B (n_0_87));
XNOR2_X1 i_0_143 (.ZN (n_0_86), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_142 (.ZN (u[53]), .A (y[53]), .B (n_0_86));
XNOR2_X1 i_0_141 (.ZN (n_0_85), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_140 (.ZN (u[52]), .A (y[52]), .B (n_0_85));
XNOR2_X1 i_0_139 (.ZN (n_0_84), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_138 (.ZN (u[51]), .A (y[51]), .B (n_0_84));
XNOR2_X1 i_0_137 (.ZN (n_0_83), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_136 (.ZN (u[50]), .A (y[50]), .B (n_0_83));
XNOR2_X1 i_0_135 (.ZN (n_0_82), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_134 (.ZN (u[49]), .A (y[49]), .B (n_0_82));
XNOR2_X1 i_0_133 (.ZN (n_0_81), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_132 (.ZN (u[48]), .A (y[48]), .B (n_0_81));
XNOR2_X1 i_0_131 (.ZN (n_0_80), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_130 (.ZN (u[47]), .A (y[47]), .B (n_0_80));
XNOR2_X1 i_0_129 (.ZN (n_0_79), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_128 (.ZN (u[46]), .A (y[46]), .B (n_0_79));
XNOR2_X1 i_0_127 (.ZN (n_0_78), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_126 (.ZN (u[45]), .A (y[45]), .B (n_0_78));
XNOR2_X1 i_0_125 (.ZN (n_0_77), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_124 (.ZN (u[44]), .A (y[44]), .B (n_0_77));
XNOR2_X1 i_0_123 (.ZN (n_0_76), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_122 (.ZN (u[43]), .A (y[43]), .B (n_0_76));
XNOR2_X1 i_0_121 (.ZN (n_0_75), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_120 (.ZN (u[42]), .A (y[42]), .B (n_0_75));
XNOR2_X1 i_0_119 (.ZN (n_0_74), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_118 (.ZN (u[41]), .A (y[41]), .B (n_0_74));
XNOR2_X1 i_0_117 (.ZN (n_0_73), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_116 (.ZN (u[40]), .A (y[40]), .B (n_0_73));
XNOR2_X1 i_0_115 (.ZN (n_0_72), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_114 (.ZN (u[39]), .A (y[39]), .B (n_0_72));
XNOR2_X1 i_0_113 (.ZN (n_0_71), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_112 (.ZN (u[38]), .A (y[38]), .B (n_0_71));
XNOR2_X1 i_0_111 (.ZN (n_0_70), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_110 (.ZN (u[37]), .A (y[37]), .B (n_0_70));
XNOR2_X1 i_0_109 (.ZN (n_0_69), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_108 (.ZN (u[36]), .A (y[36]), .B (n_0_69));
XNOR2_X1 i_0_107 (.ZN (n_0_68), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_106 (.ZN (u[35]), .A (y[35]), .B (n_0_68));
XNOR2_X1 i_0_105 (.ZN (n_0_67), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_104 (.ZN (u[34]), .A (y[34]), .B (n_0_67));
XNOR2_X1 i_0_103 (.ZN (n_0_66), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_102 (.ZN (u[33]), .A (y[33]), .B (n_0_66));
XNOR2_X1 i_0_101 (.ZN (n_0_65), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_100 (.ZN (u[32]), .A (y[32]), .B (n_0_65));
XNOR2_X1 i_0_99 (.ZN (n_0_64), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_98 (.ZN (u[31]), .A (y[31]), .B (n_0_64));
XOR2_X1 i_0_97 (.Z (u[30]), .A (y[30]), .B (x[30]));
NAND2_X1 i_0_96 (.ZN (n_0_63), .A1 (z[63]), .A2 (x[62]));
OAI21_X1 i_0_95 (.ZN (n_0_62), .A (y[62]), .B1 (z[63]), .B2 (x[62]));
NAND2_X1 i_0_94 (.ZN (v[63]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_93 (.ZN (n_0_61), .A1 (z[61]), .A2 (x[61]));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (y[61]), .B1 (z[61]), .B2 (x[61]));
NAND2_X1 i_0_91 (.ZN (v[62]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[60]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_88 (.ZN (v[61]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[59]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_85 (.ZN (v[60]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_82 (.ZN (v[59]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_79 (.ZN (v[58]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_76 (.ZN (v[57]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_73 (.ZN (v[56]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_70 (.ZN (v[55]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_67 (.ZN (v[54]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_64 (.ZN (v[53]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_61 (.ZN (v[52]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_58 (.ZN (v[51]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_55 (.ZN (v[50]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_52 (.ZN (v[49]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_49 (.ZN (v[48]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_46 (.ZN (v[47]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_43 (.ZN (v[46]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_40 (.ZN (v[45]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (y[43]), .A2 (z[43]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (x[43]), .B1 (z[43]), .B2 (y[43]));
NAND2_X1 i_0_37 (.ZN (v[44]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_34 (.ZN (v[43]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_31 (.ZN (v[42]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_28 (.ZN (v[41]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_25 (.ZN (v[40]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_22 (.ZN (v[39]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_19 (.ZN (v[38]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_16 (.ZN (v[37]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_13 (.ZN (v[36]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_10 (.ZN (v[35]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_7 (.ZN (v[34]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_4 (.ZN (v[33]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_1 (.ZN (v[32]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[31]), .A1 (y[30]), .A2 (x[30]));

endmodule //CSA__5_197

module CSA__5_194 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;


XNOR2_X1 i_0_168 (.ZN (n_0_99), .A (z[62]), .B (x[63]));
XNOR2_X1 i_0_167 (.ZN (u[63]), .A (y[63]), .B (n_0_99));
XNOR2_X1 i_0_166 (.ZN (n_0_98), .A (z[62]), .B (x[62]));
XNOR2_X1 i_0_165 (.ZN (u[62]), .A (y[62]), .B (n_0_98));
XNOR2_X1 i_0_164 (.ZN (n_0_97), .A (z[62]), .B (x[61]));
XNOR2_X1 i_0_163 (.ZN (u[61]), .A (y[61]), .B (n_0_97));
XNOR2_X1 i_0_162 (.ZN (n_0_96), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_161 (.ZN (u[60]), .A (y[60]), .B (n_0_96));
XNOR2_X1 i_0_160 (.ZN (n_0_95), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_159 (.ZN (u[59]), .A (y[59]), .B (n_0_95));
XNOR2_X1 i_0_158 (.ZN (n_0_94), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_157 (.ZN (u[58]), .A (y[58]), .B (n_0_94));
XNOR2_X1 i_0_156 (.ZN (n_0_93), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_155 (.ZN (u[57]), .A (y[57]), .B (n_0_93));
XNOR2_X1 i_0_154 (.ZN (n_0_92), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_153 (.ZN (u[56]), .A (y[56]), .B (n_0_92));
XNOR2_X1 i_0_152 (.ZN (n_0_91), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_151 (.ZN (u[55]), .A (y[55]), .B (n_0_91));
XNOR2_X1 i_0_150 (.ZN (n_0_90), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_149 (.ZN (u[54]), .A (y[54]), .B (n_0_90));
XNOR2_X1 i_0_148 (.ZN (n_0_89), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_147 (.ZN (u[53]), .A (y[53]), .B (n_0_89));
XNOR2_X1 i_0_146 (.ZN (n_0_88), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_145 (.ZN (u[52]), .A (y[52]), .B (n_0_88));
XNOR2_X1 i_0_144 (.ZN (n_0_87), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_143 (.ZN (u[51]), .A (y[51]), .B (n_0_87));
XNOR2_X1 i_0_142 (.ZN (n_0_86), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_141 (.ZN (u[50]), .A (y[50]), .B (n_0_86));
XNOR2_X1 i_0_140 (.ZN (n_0_85), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_139 (.ZN (u[49]), .A (y[49]), .B (n_0_85));
XNOR2_X1 i_0_138 (.ZN (n_0_84), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_137 (.ZN (u[48]), .A (y[48]), .B (n_0_84));
XNOR2_X1 i_0_136 (.ZN (n_0_83), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_135 (.ZN (u[47]), .A (y[47]), .B (n_0_83));
XNOR2_X1 i_0_134 (.ZN (n_0_82), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_133 (.ZN (u[46]), .A (y[46]), .B (n_0_82));
XNOR2_X1 i_0_132 (.ZN (n_0_81), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_131 (.ZN (u[45]), .A (y[45]), .B (n_0_81));
XNOR2_X1 i_0_130 (.ZN (n_0_80), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_129 (.ZN (u[44]), .A (y[44]), .B (n_0_80));
XNOR2_X1 i_0_128 (.ZN (n_0_79), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_127 (.ZN (u[43]), .A (y[43]), .B (n_0_79));
XNOR2_X1 i_0_126 (.ZN (n_0_78), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_125 (.ZN (u[42]), .A (y[42]), .B (n_0_78));
XNOR2_X1 i_0_124 (.ZN (n_0_77), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_123 (.ZN (u[41]), .A (y[41]), .B (n_0_77));
XNOR2_X1 i_0_122 (.ZN (n_0_76), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_121 (.ZN (u[40]), .A (y[40]), .B (n_0_76));
XNOR2_X1 i_0_120 (.ZN (n_0_75), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_119 (.ZN (u[39]), .A (y[39]), .B (n_0_75));
XNOR2_X1 i_0_118 (.ZN (n_0_74), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_117 (.ZN (u[38]), .A (y[38]), .B (n_0_74));
XNOR2_X1 i_0_116 (.ZN (n_0_73), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_115 (.ZN (u[37]), .A (y[37]), .B (n_0_73));
XNOR2_X1 i_0_114 (.ZN (n_0_72), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_113 (.ZN (u[36]), .A (y[36]), .B (n_0_72));
XNOR2_X1 i_0_112 (.ZN (n_0_71), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_111 (.ZN (u[35]), .A (y[35]), .B (n_0_71));
XNOR2_X1 i_0_110 (.ZN (n_0_70), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_109 (.ZN (u[34]), .A (y[34]), .B (n_0_70));
XNOR2_X1 i_0_108 (.ZN (n_0_69), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_107 (.ZN (u[33]), .A (y[33]), .B (n_0_69));
XNOR2_X1 i_0_106 (.ZN (n_0_68), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_105 (.ZN (u[32]), .A (y[32]), .B (n_0_68));
XNOR2_X1 i_0_104 (.ZN (n_0_67), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_103 (.ZN (u[31]), .A (y[31]), .B (n_0_67));
XNOR2_X1 i_0_102 (.ZN (n_0_66), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_101 (.ZN (u[30]), .A (y[30]), .B (n_0_66));
XOR2_X1 i_0_100 (.Z (u[29]), .A (y[29]), .B (x[29]));
NAND2_X1 i_0_99 (.ZN (n_0_65), .A1 (z[62]), .A2 (x[62]));
OAI21_X1 i_0_98 (.ZN (n_0_64), .A (y[62]), .B1 (z[62]), .B2 (x[62]));
NAND2_X1 i_0_97 (.ZN (v[63]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_96 (.ZN (n_0_63), .A1 (z[62]), .A2 (x[61]));
OAI21_X1 i_0_95 (.ZN (n_0_62), .A (y[61]), .B1 (z[62]), .B2 (x[61]));
NAND2_X1 i_0_94 (.ZN (v[62]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_93 (.ZN (n_0_61), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (y[60]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_91 (.ZN (v[61]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[59]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_88 (.ZN (v[60]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_85 (.ZN (v[59]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_82 (.ZN (v[58]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_79 (.ZN (v[57]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_76 (.ZN (v[56]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_73 (.ZN (v[55]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_70 (.ZN (v[54]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_67 (.ZN (v[53]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_64 (.ZN (v[52]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_61 (.ZN (v[51]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_58 (.ZN (v[50]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_55 (.ZN (v[49]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_52 (.ZN (v[48]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_49 (.ZN (v[47]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (y[45]), .A2 (z[45]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (x[45]), .B1 (z[45]), .B2 (y[45]));
NAND2_X1 i_0_46 (.ZN (v[46]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_43 (.ZN (v[45]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_40 (.ZN (v[44]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_37 (.ZN (v[43]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_34 (.ZN (v[42]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_31 (.ZN (v[41]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_28 (.ZN (v[40]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_25 (.ZN (v[39]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_22 (.ZN (v[38]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_19 (.ZN (v[37]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_16 (.ZN (v[36]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_13 (.ZN (v[35]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_10 (.ZN (v[34]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_7 (.ZN (v[33]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_4 (.ZN (v[32]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_1 (.ZN (v[31]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[30]), .A1 (y[29]), .A2 (x[29]));

endmodule //CSA__5_194

module CSA__5_191 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;


INV_X1 i_0_169 (.ZN (n_0_98), .A (x[62]));
INV_X1 i_0_168 (.ZN (n_0_97), .A (x[61]));
INV_X1 i_0_167 (.ZN (n_0_96), .A (x[60]));
XOR2_X1 i_0_166 (.Z (n_0_95), .A (y[62]), .B (z[62]));
XOR2_X1 i_0_165 (.Z (u[63]), .A (x[63]), .B (n_0_95));
XNOR2_X1 i_0_164 (.ZN (u[62]), .A (n_0_98), .B (n_0_95));
XNOR2_X1 i_0_163 (.ZN (u[61]), .A (n_0_97), .B (n_0_95));
XNOR2_X1 i_0_162 (.ZN (u[60]), .A (n_0_96), .B (n_0_95));
XNOR2_X1 i_0_161 (.ZN (n_0_94), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_160 (.ZN (u[59]), .A (y[62]), .B (n_0_94));
XNOR2_X1 i_0_159 (.ZN (n_0_93), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_158 (.ZN (u[58]), .A (y[58]), .B (n_0_93));
XNOR2_X1 i_0_157 (.ZN (n_0_92), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_156 (.ZN (u[57]), .A (y[57]), .B (n_0_92));
XNOR2_X1 i_0_155 (.ZN (n_0_91), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_154 (.ZN (u[56]), .A (y[56]), .B (n_0_91));
XNOR2_X1 i_0_153 (.ZN (n_0_90), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_152 (.ZN (u[55]), .A (y[55]), .B (n_0_90));
XNOR2_X1 i_0_151 (.ZN (n_0_89), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_150 (.ZN (u[54]), .A (y[54]), .B (n_0_89));
XNOR2_X1 i_0_149 (.ZN (n_0_88), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_148 (.ZN (u[53]), .A (y[53]), .B (n_0_88));
XNOR2_X1 i_0_147 (.ZN (n_0_87), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_146 (.ZN (u[52]), .A (y[52]), .B (n_0_87));
XNOR2_X1 i_0_145 (.ZN (n_0_86), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_144 (.ZN (u[51]), .A (y[51]), .B (n_0_86));
XNOR2_X1 i_0_143 (.ZN (n_0_85), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_142 (.ZN (u[50]), .A (y[50]), .B (n_0_85));
XNOR2_X1 i_0_141 (.ZN (n_0_84), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_140 (.ZN (u[49]), .A (y[49]), .B (n_0_84));
XNOR2_X1 i_0_139 (.ZN (n_0_83), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_138 (.ZN (u[48]), .A (y[48]), .B (n_0_83));
XNOR2_X1 i_0_137 (.ZN (n_0_82), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_136 (.ZN (u[47]), .A (y[47]), .B (n_0_82));
XNOR2_X1 i_0_135 (.ZN (n_0_81), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_134 (.ZN (u[46]), .A (y[46]), .B (n_0_81));
XNOR2_X1 i_0_133 (.ZN (n_0_80), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_132 (.ZN (u[45]), .A (y[45]), .B (n_0_80));
XNOR2_X1 i_0_131 (.ZN (n_0_79), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_130 (.ZN (u[44]), .A (y[44]), .B (n_0_79));
XNOR2_X1 i_0_129 (.ZN (n_0_78), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_128 (.ZN (u[43]), .A (y[43]), .B (n_0_78));
XNOR2_X1 i_0_127 (.ZN (n_0_77), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_126 (.ZN (u[42]), .A (y[42]), .B (n_0_77));
XNOR2_X1 i_0_125 (.ZN (n_0_76), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_124 (.ZN (u[41]), .A (y[41]), .B (n_0_76));
XNOR2_X1 i_0_123 (.ZN (n_0_75), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_122 (.ZN (u[40]), .A (y[40]), .B (n_0_75));
XNOR2_X1 i_0_121 (.ZN (n_0_74), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_120 (.ZN (u[39]), .A (y[39]), .B (n_0_74));
XNOR2_X1 i_0_119 (.ZN (n_0_73), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_118 (.ZN (u[38]), .A (y[38]), .B (n_0_73));
XNOR2_X1 i_0_117 (.ZN (n_0_72), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_116 (.ZN (u[37]), .A (y[37]), .B (n_0_72));
XNOR2_X1 i_0_115 (.ZN (n_0_71), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_114 (.ZN (u[36]), .A (y[36]), .B (n_0_71));
XNOR2_X1 i_0_113 (.ZN (n_0_70), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_112 (.ZN (u[35]), .A (y[35]), .B (n_0_70));
XNOR2_X1 i_0_111 (.ZN (n_0_69), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_110 (.ZN (u[34]), .A (y[34]), .B (n_0_69));
XNOR2_X1 i_0_109 (.ZN (n_0_68), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_108 (.ZN (u[33]), .A (y[33]), .B (n_0_68));
XNOR2_X1 i_0_107 (.ZN (n_0_67), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_106 (.ZN (u[32]), .A (y[32]), .B (n_0_67));
XNOR2_X1 i_0_105 (.ZN (n_0_66), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_104 (.ZN (u[31]), .A (y[31]), .B (n_0_66));
XNOR2_X1 i_0_103 (.ZN (n_0_65), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_102 (.ZN (u[30]), .A (y[30]), .B (n_0_65));
XNOR2_X1 i_0_101 (.ZN (n_0_64), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_100 (.ZN (u[29]), .A (y[29]), .B (n_0_64));
XOR2_X1 i_0_99 (.Z (u[28]), .A (y[28]), .B (x[28]));
NAND2_X1 i_0_98 (.ZN (n_0_63), .A1 (y[62]), .A2 (z[62]));
NOR2_X1 i_0_97 (.ZN (n_0_62), .A1 (y[62]), .A2 (z[62]));
OAI21_X1 i_0_96 (.ZN (v[63]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_98));
OAI21_X1 i_0_95 (.ZN (v[62]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_97));
OAI21_X1 i_0_94 (.ZN (v[61]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_96));
NAND2_X1 i_0_93 (.ZN (n_0_61), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (y[62]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_91 (.ZN (v[60]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_88 (.ZN (v[59]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_85 (.ZN (v[58]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_82 (.ZN (v[57]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_79 (.ZN (v[56]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_76 (.ZN (v[55]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_73 (.ZN (v[54]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_70 (.ZN (v[53]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_67 (.ZN (v[52]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_64 (.ZN (v[51]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_61 (.ZN (v[50]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_58 (.ZN (v[49]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_55 (.ZN (v[48]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_52 (.ZN (v[47]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_49 (.ZN (v[46]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_46 (.ZN (v[45]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_43 (.ZN (v[44]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_40 (.ZN (v[43]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_37 (.ZN (v[42]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_34 (.ZN (v[41]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_31 (.ZN (v[40]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_28 (.ZN (v[39]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_25 (.ZN (v[38]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_22 (.ZN (v[37]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_19 (.ZN (v[36]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_16 (.ZN (v[35]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_13 (.ZN (v[34]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_10 (.ZN (v[33]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_7 (.ZN (v[32]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_4 (.ZN (v[31]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_1 (.ZN (v[30]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[29]), .A1 (y[28]), .A2 (x[28]));

endmodule //CSA__5_191

module CSA__0_78 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;


XOR2_X1 i_0_176 (.Z (n_0_102), .A (y[63]), .B (x[63]));
XOR2_X2 i_0_175 (.Z (u[63]), .A (z[63]), .B (n_0_102));
XOR2_X1 i_0_174 (.Z (u[58]), .A (z[58]), .B (n_0_102));
XNOR2_X1 i_0_173 (.ZN (n_0_101), .A (z[57]), .B (x[63]));
XNOR2_X1 i_0_172 (.ZN (u[57]), .A (y[57]), .B (n_0_101));
XNOR2_X1 i_0_171 (.ZN (n_0_100), .A (z[56]), .B (x[63]));
XNOR2_X1 i_0_170 (.ZN (u[56]), .A (y[56]), .B (n_0_100));
XNOR2_X1 i_0_169 (.ZN (n_0_99), .A (z[55]), .B (x[63]));
XNOR2_X1 i_0_168 (.ZN (u[55]), .A (y[55]), .B (n_0_99));
XNOR2_X1 i_0_167 (.ZN (n_0_98), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_166 (.ZN (u[54]), .A (y[54]), .B (n_0_98));
XNOR2_X1 i_0_165 (.ZN (n_0_97), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_164 (.ZN (u[53]), .A (y[53]), .B (n_0_97));
XNOR2_X1 i_0_163 (.ZN (n_0_96), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_162 (.ZN (u[52]), .A (y[52]), .B (n_0_96));
XNOR2_X1 i_0_161 (.ZN (n_0_95), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_160 (.ZN (u[51]), .A (y[51]), .B (n_0_95));
XNOR2_X1 i_0_159 (.ZN (n_0_94), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_158 (.ZN (u[50]), .A (y[50]), .B (n_0_94));
XNOR2_X1 i_0_157 (.ZN (n_0_93), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_156 (.ZN (u[49]), .A (y[49]), .B (n_0_93));
XNOR2_X1 i_0_155 (.ZN (n_0_92), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_154 (.ZN (u[48]), .A (y[48]), .B (n_0_92));
XNOR2_X1 i_0_153 (.ZN (n_0_91), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_152 (.ZN (u[47]), .A (y[47]), .B (n_0_91));
XNOR2_X1 i_0_151 (.ZN (n_0_90), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_150 (.ZN (u[46]), .A (y[46]), .B (n_0_90));
XNOR2_X1 i_0_149 (.ZN (n_0_89), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_148 (.ZN (u[45]), .A (y[45]), .B (n_0_89));
XNOR2_X1 i_0_147 (.ZN (n_0_88), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_146 (.ZN (u[44]), .A (y[44]), .B (n_0_88));
XNOR2_X1 i_0_145 (.ZN (n_0_87), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_144 (.ZN (u[43]), .A (y[43]), .B (n_0_87));
XNOR2_X1 i_0_143 (.ZN (n_0_86), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_142 (.ZN (u[42]), .A (y[42]), .B (n_0_86));
XNOR2_X1 i_0_141 (.ZN (n_0_85), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_140 (.ZN (u[41]), .A (y[41]), .B (n_0_85));
XNOR2_X1 i_0_139 (.ZN (n_0_84), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_138 (.ZN (u[40]), .A (y[40]), .B (n_0_84));
XNOR2_X1 i_0_137 (.ZN (n_0_83), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_136 (.ZN (u[39]), .A (y[39]), .B (n_0_83));
XNOR2_X1 i_0_135 (.ZN (n_0_82), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_134 (.ZN (u[38]), .A (y[38]), .B (n_0_82));
XNOR2_X1 i_0_133 (.ZN (n_0_81), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_132 (.ZN (u[37]), .A (y[37]), .B (n_0_81));
XNOR2_X1 i_0_131 (.ZN (n_0_80), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_130 (.ZN (u[36]), .A (y[36]), .B (n_0_80));
XNOR2_X1 i_0_129 (.ZN (n_0_79), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_128 (.ZN (u[35]), .A (y[35]), .B (n_0_79));
XNOR2_X1 i_0_127 (.ZN (n_0_78), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_126 (.ZN (u[34]), .A (y[34]), .B (n_0_78));
XNOR2_X1 i_0_125 (.ZN (n_0_77), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_124 (.ZN (u[33]), .A (y[33]), .B (n_0_77));
XNOR2_X1 i_0_123 (.ZN (n_0_76), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_122 (.ZN (u[32]), .A (y[32]), .B (n_0_76));
XNOR2_X1 i_0_121 (.ZN (n_0_75), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_120 (.ZN (u[31]), .A (y[31]), .B (n_0_75));
XNOR2_X1 i_0_119 (.ZN (n_0_74), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_118 (.ZN (u[30]), .A (y[30]), .B (n_0_74));
XNOR2_X1 i_0_117 (.ZN (n_0_73), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_116 (.ZN (u[29]), .A (y[29]), .B (n_0_73));
XNOR2_X1 i_0_115 (.ZN (n_0_72), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_114 (.ZN (u[28]), .A (y[28]), .B (n_0_72));
XNOR2_X1 i_0_113 (.ZN (n_0_71), .A (z[27]), .B (x[27]));
XNOR2_X2 i_0_112 (.ZN (u[27]), .A (y[27]), .B (n_0_71));
XNOR2_X1 i_0_111 (.ZN (n_0_70), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_110 (.ZN (u[26]), .A (y[26]), .B (n_0_70));
XNOR2_X1 i_0_109 (.ZN (n_0_69), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_108 (.ZN (u[25]), .A (y[25]), .B (n_0_69));
XOR2_X1 i_0_107 (.Z (u[24]), .A (y[24]), .B (x[24]));
XOR2_X1 i_0_106 (.Z (u[23]), .A (y[23]), .B (x[23]));
NAND2_X1 i_0_105 (.ZN (n_0_68), .A1 (y[63]), .A2 (x[63]));
OAI21_X1 i_0_104 (.ZN (n_0_67), .A (z[63]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_103 (.ZN (v[63]), .A1 (n_0_68), .A2 (n_0_67));
OAI21_X1 i_0_102 (.ZN (n_0_66), .A (z[58]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_101 (.ZN (v[59]), .A1 (n_0_68), .A2 (n_0_66));
NAND2_X1 i_0_100 (.ZN (n_0_65), .A1 (z[57]), .A2 (x[63]));
OAI21_X1 i_0_99 (.ZN (n_0_64), .A (y[57]), .B1 (z[57]), .B2 (x[63]));
NAND2_X1 i_0_98 (.ZN (v[58]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_97 (.ZN (n_0_63), .A1 (z[56]), .A2 (x[63]));
OAI21_X1 i_0_96 (.ZN (n_0_62), .A (y[56]), .B1 (z[56]), .B2 (x[63]));
NAND2_X1 i_0_95 (.ZN (v[57]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_94 (.ZN (n_0_61), .A1 (z[55]), .A2 (x[63]));
OAI21_X1 i_0_93 (.ZN (n_0_60), .A (y[55]), .B1 (z[55]), .B2 (x[63]));
NAND2_X1 i_0_92 (.ZN (v[56]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_91 (.ZN (n_0_59), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_90 (.ZN (n_0_58), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_89 (.ZN (v[55]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_88 (.ZN (n_0_57), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_87 (.ZN (n_0_56), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_86 (.ZN (v[54]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_85 (.ZN (n_0_55), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_84 (.ZN (n_0_54), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_83 (.ZN (v[53]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_82 (.ZN (n_0_53), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_81 (.ZN (n_0_52), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_80 (.ZN (v[52]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_79 (.ZN (n_0_51), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_78 (.ZN (n_0_50), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_77 (.ZN (v[51]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_76 (.ZN (n_0_49), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_75 (.ZN (n_0_48), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_74 (.ZN (v[50]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_73 (.ZN (n_0_47), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_72 (.ZN (n_0_46), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_71 (.ZN (v[49]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_70 (.ZN (n_0_45), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_69 (.ZN (n_0_44), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_68 (.ZN (v[48]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_67 (.ZN (n_0_43), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_66 (.ZN (n_0_42), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_65 (.ZN (v[47]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_64 (.ZN (n_0_41), .A1 (y[45]), .A2 (z[45]));
OAI21_X1 i_0_63 (.ZN (n_0_40), .A (x[45]), .B1 (z[45]), .B2 (y[45]));
NAND2_X1 i_0_62 (.ZN (v[46]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_61 (.ZN (n_0_39), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_60 (.ZN (n_0_38), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_59 (.ZN (v[45]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_58 (.ZN (n_0_37), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_57 (.ZN (n_0_36), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_56 (.ZN (v[44]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_55 (.ZN (n_0_35), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_54 (.ZN (n_0_34), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_53 (.ZN (v[43]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_52 (.ZN (n_0_33), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_51 (.ZN (n_0_32), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_50 (.ZN (v[42]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_49 (.ZN (n_0_31), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_48 (.ZN (n_0_30), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_47 (.ZN (v[41]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_46 (.ZN (n_0_29), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_45 (.ZN (n_0_28), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_44 (.ZN (v[40]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_43 (.ZN (n_0_27), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_42 (.ZN (n_0_26), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_41 (.ZN (v[39]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_40 (.ZN (n_0_25), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_39 (.ZN (n_0_24), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_38 (.ZN (v[38]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_37 (.ZN (n_0_23), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_36 (.ZN (n_0_22), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_35 (.ZN (v[37]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_34 (.ZN (n_0_21), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_33 (.ZN (n_0_20), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_32 (.ZN (v[36]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_31 (.ZN (n_0_19), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_30 (.ZN (n_0_18), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_29 (.ZN (v[35]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_28 (.ZN (n_0_17), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_27 (.ZN (n_0_16), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_26 (.ZN (v[34]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_25 (.ZN (n_0_15), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_24 (.ZN (n_0_14), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_23 (.ZN (v[33]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_22 (.ZN (n_0_13), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_21 (.ZN (n_0_12), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_20 (.ZN (v[32]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_19 (.ZN (n_0_11), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_18 (.ZN (n_0_10), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_17 (.ZN (v[31]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_16 (.ZN (n_0_9), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_15 (.ZN (n_0_8), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_14 (.ZN (v[30]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_13 (.ZN (n_0_7), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_12 (.ZN (n_0_6), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_11 (.ZN (v[29]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_10 (.ZN (n_0_5), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_9 (.ZN (n_0_4), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_8 (.ZN (v[28]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_7 (.ZN (n_0_3), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_6 (.ZN (n_0_2), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_5 (.ZN (v[27]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_4 (.ZN (n_0_1), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_3 (.ZN (n_0_0), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_2 (.ZN (v[26]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_1 (.ZN (v[25]), .A1 (y[24]), .A2 (x[24]));
AND2_X1 i_0_0 (.ZN (v[24]), .A1 (y[23]), .A2 (x[23]));

endmodule //CSA__0_78

module CSA__4_20 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;


XOR2_X1 i_0_166 (.Z (n_0_96), .A (y[63]), .B (x[63]));
XOR2_X1 i_0_165 (.Z (u[63]), .A (z[63]), .B (n_0_96));
XOR2_X1 i_0_164 (.Z (u[57]), .A (z[57]), .B (n_0_96));
XNOR2_X1 i_0_163 (.ZN (n_0_95), .A (z[56]), .B (x[63]));
XNOR2_X1 i_0_162 (.ZN (u[56]), .A (y[56]), .B (n_0_95));
XNOR2_X1 i_0_161 (.ZN (n_0_94), .A (z[55]), .B (x[63]));
XNOR2_X1 i_0_160 (.ZN (u[55]), .A (y[55]), .B (n_0_94));
XNOR2_X1 i_0_159 (.ZN (n_0_93), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_158 (.ZN (u[54]), .A (y[54]), .B (n_0_93));
XNOR2_X1 i_0_157 (.ZN (n_0_92), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_156 (.ZN (u[53]), .A (y[53]), .B (n_0_92));
XNOR2_X1 i_0_155 (.ZN (n_0_91), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_154 (.ZN (u[52]), .A (y[52]), .B (n_0_91));
XNOR2_X1 i_0_153 (.ZN (n_0_90), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_152 (.ZN (u[51]), .A (y[51]), .B (n_0_90));
XNOR2_X1 i_0_151 (.ZN (n_0_89), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_150 (.ZN (u[50]), .A (y[50]), .B (n_0_89));
XNOR2_X1 i_0_149 (.ZN (n_0_88), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_148 (.ZN (u[49]), .A (y[49]), .B (n_0_88));
XNOR2_X1 i_0_147 (.ZN (n_0_87), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_146 (.ZN (u[48]), .A (y[48]), .B (n_0_87));
XNOR2_X1 i_0_145 (.ZN (n_0_86), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_144 (.ZN (u[47]), .A (y[47]), .B (n_0_86));
XNOR2_X1 i_0_143 (.ZN (n_0_85), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_142 (.ZN (u[46]), .A (y[46]), .B (n_0_85));
XNOR2_X1 i_0_141 (.ZN (n_0_84), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_140 (.ZN (u[45]), .A (y[45]), .B (n_0_84));
XNOR2_X1 i_0_139 (.ZN (n_0_83), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_138 (.ZN (u[44]), .A (y[44]), .B (n_0_83));
XNOR2_X1 i_0_137 (.ZN (n_0_82), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_136 (.ZN (u[43]), .A (y[43]), .B (n_0_82));
XNOR2_X1 i_0_135 (.ZN (n_0_81), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_134 (.ZN (u[42]), .A (y[42]), .B (n_0_81));
XNOR2_X1 i_0_133 (.ZN (n_0_80), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_132 (.ZN (u[41]), .A (y[41]), .B (n_0_80));
XNOR2_X1 i_0_131 (.ZN (n_0_79), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_130 (.ZN (u[40]), .A (y[40]), .B (n_0_79));
XNOR2_X1 i_0_129 (.ZN (n_0_78), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_128 (.ZN (u[39]), .A (y[39]), .B (n_0_78));
XNOR2_X1 i_0_127 (.ZN (n_0_77), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_126 (.ZN (u[38]), .A (y[38]), .B (n_0_77));
XNOR2_X1 i_0_125 (.ZN (n_0_76), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_124 (.ZN (u[37]), .A (y[37]), .B (n_0_76));
XNOR2_X1 i_0_123 (.ZN (n_0_75), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_122 (.ZN (u[36]), .A (y[36]), .B (n_0_75));
XNOR2_X1 i_0_121 (.ZN (n_0_74), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_120 (.ZN (u[35]), .A (y[35]), .B (n_0_74));
XNOR2_X1 i_0_119 (.ZN (n_0_73), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_118 (.ZN (u[34]), .A (y[34]), .B (n_0_73));
XNOR2_X1 i_0_117 (.ZN (n_0_72), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_116 (.ZN (u[33]), .A (y[33]), .B (n_0_72));
XNOR2_X1 i_0_115 (.ZN (n_0_71), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_114 (.ZN (u[32]), .A (y[32]), .B (n_0_71));
XNOR2_X1 i_0_113 (.ZN (n_0_70), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_112 (.ZN (u[31]), .A (y[31]), .B (n_0_70));
XNOR2_X1 i_0_111 (.ZN (n_0_69), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_110 (.ZN (u[30]), .A (y[30]), .B (n_0_69));
XNOR2_X1 i_0_109 (.ZN (n_0_68), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_108 (.ZN (u[29]), .A (y[29]), .B (n_0_68));
XNOR2_X1 i_0_107 (.ZN (n_0_67), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_106 (.ZN (u[28]), .A (y[28]), .B (n_0_67));
XNOR2_X1 i_0_105 (.ZN (n_0_66), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_104 (.ZN (u[27]), .A (y[27]), .B (n_0_66));
XNOR2_X1 i_0_103 (.ZN (n_0_65), .A (z[26]), .B (x[26]));
XNOR2_X2 i_0_102 (.ZN (u[26]), .A (y[26]), .B (n_0_65));
XOR2_X1 i_0_101 (.Z (u[25]), .A (y[25]), .B (x[25]));
XOR2_X1 i_0_100 (.Z (u[24]), .A (y[24]), .B (x[24]));
NAND2_X1 i_0_99 (.ZN (n_0_64), .A1 (y[63]), .A2 (x[63]));
OAI21_X1 i_0_98 (.ZN (n_0_63), .A (z[63]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_97 (.ZN (v[63]), .A1 (n_0_64), .A2 (n_0_63));
OAI21_X1 i_0_96 (.ZN (n_0_62), .A (z[57]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_95 (.ZN (v[58]), .A1 (n_0_64), .A2 (n_0_62));
NAND2_X1 i_0_94 (.ZN (n_0_61), .A1 (z[56]), .A2 (x[63]));
OAI21_X1 i_0_93 (.ZN (n_0_60), .A (y[56]), .B1 (z[56]), .B2 (x[63]));
NAND2_X1 i_0_92 (.ZN (v[57]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_91 (.ZN (n_0_59), .A1 (z[55]), .A2 (x[63]));
OAI21_X1 i_0_90 (.ZN (n_0_58), .A (y[55]), .B1 (z[55]), .B2 (x[63]));
NAND2_X1 i_0_89 (.ZN (v[56]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_88 (.ZN (n_0_57), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_87 (.ZN (n_0_56), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_86 (.ZN (v[55]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_85 (.ZN (n_0_55), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_84 (.ZN (n_0_54), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_83 (.ZN (v[54]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_82 (.ZN (n_0_53), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_81 (.ZN (n_0_52), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_80 (.ZN (v[53]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_79 (.ZN (n_0_51), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_78 (.ZN (n_0_50), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_77 (.ZN (v[52]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_76 (.ZN (n_0_49), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_75 (.ZN (n_0_48), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_74 (.ZN (v[51]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_73 (.ZN (n_0_47), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_72 (.ZN (n_0_46), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_71 (.ZN (v[50]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_70 (.ZN (n_0_45), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_69 (.ZN (n_0_44), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_68 (.ZN (v[49]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_67 (.ZN (n_0_43), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_66 (.ZN (n_0_42), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_65 (.ZN (v[48]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_64 (.ZN (n_0_41), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_63 (.ZN (n_0_40), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_62 (.ZN (v[47]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_61 (.ZN (n_0_39), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_60 (.ZN (n_0_38), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_59 (.ZN (v[46]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_58 (.ZN (n_0_37), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_57 (.ZN (n_0_36), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_56 (.ZN (v[45]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_55 (.ZN (n_0_35), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_54 (.ZN (n_0_34), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_53 (.ZN (v[44]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_52 (.ZN (n_0_33), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_51 (.ZN (n_0_32), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_50 (.ZN (v[43]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_49 (.ZN (n_0_31), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_48 (.ZN (n_0_30), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_47 (.ZN (v[42]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_46 (.ZN (n_0_29), .A1 (y[40]), .A2 (z[40]));
OAI21_X1 i_0_45 (.ZN (n_0_28), .A (x[40]), .B1 (z[40]), .B2 (y[40]));
NAND2_X1 i_0_44 (.ZN (v[41]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_43 (.ZN (n_0_27), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_42 (.ZN (n_0_26), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_41 (.ZN (v[40]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_40 (.ZN (n_0_25), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_39 (.ZN (n_0_24), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_38 (.ZN (v[39]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_37 (.ZN (n_0_23), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_36 (.ZN (n_0_22), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_35 (.ZN (v[38]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_34 (.ZN (n_0_21), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_33 (.ZN (n_0_20), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_32 (.ZN (v[37]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_31 (.ZN (n_0_19), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_30 (.ZN (n_0_18), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_29 (.ZN (v[36]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_28 (.ZN (n_0_17), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_27 (.ZN (n_0_16), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_26 (.ZN (v[35]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_25 (.ZN (n_0_15), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_24 (.ZN (n_0_14), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_23 (.ZN (v[34]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_22 (.ZN (n_0_13), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_21 (.ZN (n_0_12), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_20 (.ZN (v[33]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_19 (.ZN (n_0_11), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_18 (.ZN (n_0_10), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_17 (.ZN (v[32]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_16 (.ZN (n_0_9), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_15 (.ZN (n_0_8), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_14 (.ZN (v[31]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_13 (.ZN (n_0_7), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_12 (.ZN (n_0_6), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_11 (.ZN (v[30]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_10 (.ZN (n_0_5), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_9 (.ZN (n_0_4), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_8 (.ZN (v[29]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_7 (.ZN (n_0_3), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_6 (.ZN (n_0_2), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_5 (.ZN (v[28]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_4 (.ZN (n_0_1), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_3 (.ZN (n_0_0), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_2 (.ZN (v[27]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_1 (.ZN (v[26]), .A1 (y[25]), .A2 (x[25]));
AND2_X1 i_0_0 (.ZN (v[25]), .A1 (y[24]), .A2 (x[24]));

endmodule //CSA__4_20

module CSA__4_17 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;


XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[63]), .B (x[63]));
XOR2_X1 i_0_158 (.Z (u[63]), .A (z[63]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[56]), .A (z[56]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[55]), .B (x[63]));
XNOR2_X1 i_0_155 (.ZN (u[55]), .A (y[55]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_153 (.ZN (u[54]), .A (y[54]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_151 (.ZN (u[53]), .A (y[53]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_149 (.ZN (u[52]), .A (y[52]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_147 (.ZN (u[51]), .A (y[51]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_145 (.ZN (u[50]), .A (y[50]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_143 (.ZN (u[49]), .A (y[49]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_141 (.ZN (u[48]), .A (y[48]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_139 (.ZN (u[47]), .A (y[47]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_137 (.ZN (u[46]), .A (y[46]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_135 (.ZN (u[45]), .A (y[45]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_133 (.ZN (u[44]), .A (y[44]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_131 (.ZN (u[43]), .A (y[43]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_129 (.ZN (u[42]), .A (y[42]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_127 (.ZN (u[41]), .A (y[41]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_125 (.ZN (u[40]), .A (y[40]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_123 (.ZN (u[39]), .A (y[39]), .B (n_0_76));
XNOR2_X1 i_0_122 (.ZN (n_0_75), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_121 (.ZN (u[38]), .A (y[38]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_119 (.ZN (u[37]), .A (y[37]), .B (n_0_74));
XNOR2_X1 i_0_118 (.ZN (n_0_73), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_117 (.ZN (u[36]), .A (y[36]), .B (n_0_73));
XNOR2_X1 i_0_116 (.ZN (n_0_72), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_115 (.ZN (u[35]), .A (y[35]), .B (n_0_72));
XNOR2_X1 i_0_114 (.ZN (n_0_71), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_113 (.ZN (u[34]), .A (y[34]), .B (n_0_71));
XNOR2_X1 i_0_112 (.ZN (n_0_70), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_111 (.ZN (u[33]), .A (y[33]), .B (n_0_70));
XNOR2_X1 i_0_110 (.ZN (n_0_69), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_109 (.ZN (u[32]), .A (y[32]), .B (n_0_69));
XNOR2_X1 i_0_108 (.ZN (n_0_68), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_107 (.ZN (u[31]), .A (y[31]), .B (n_0_68));
XNOR2_X1 i_0_106 (.ZN (n_0_67), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_105 (.ZN (u[30]), .A (y[30]), .B (n_0_67));
XNOR2_X1 i_0_104 (.ZN (n_0_66), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_103 (.ZN (u[29]), .A (y[29]), .B (n_0_66));
XNOR2_X1 i_0_102 (.ZN (n_0_65), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_101 (.ZN (u[28]), .A (y[28]), .B (n_0_65));
XNOR2_X1 i_0_100 (.ZN (n_0_64), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_99 (.ZN (u[27]), .A (y[27]), .B (n_0_64));
XNOR2_X1 i_0_98 (.ZN (n_0_63), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_97 (.ZN (u[26]), .A (y[26]), .B (n_0_63));
XOR2_X1 i_0_96 (.Z (u[25]), .A (y[25]), .B (x[25]));
NAND2_X1 i_0_95 (.ZN (n_0_62), .A1 (y[63]), .A2 (x[63]));
OAI21_X1 i_0_94 (.ZN (n_0_61), .A (z[63]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_93 (.ZN (v[63]), .A1 (n_0_62), .A2 (n_0_61));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (z[56]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_91 (.ZN (v[57]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[55]), .A2 (x[63]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[55]), .B1 (z[55]), .B2 (x[63]));
NAND2_X1 i_0_88 (.ZN (v[56]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_85 (.ZN (v[55]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_82 (.ZN (v[54]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_79 (.ZN (v[53]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_76 (.ZN (v[52]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_73 (.ZN (v[51]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_70 (.ZN (v[50]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_67 (.ZN (v[49]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_64 (.ZN (v[48]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_61 (.ZN (v[47]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_58 (.ZN (v[46]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_55 (.ZN (v[45]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_52 (.ZN (v[44]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_49 (.ZN (v[43]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_46 (.ZN (v[42]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_43 (.ZN (v[41]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_40 (.ZN (v[40]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_37 (.ZN (v[39]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_34 (.ZN (v[38]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_31 (.ZN (v[37]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_28 (.ZN (v[36]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_25 (.ZN (v[35]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_22 (.ZN (v[34]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_19 (.ZN (v[33]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_16 (.ZN (v[32]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_13 (.ZN (v[31]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_10 (.ZN (v[30]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_7 (.ZN (v[29]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_4 (.ZN (v[28]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_1 (.ZN (v[27]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[26]), .A1 (y[25]), .A2 (x[25]));

endmodule //CSA__4_17

module CSA__4_14 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;


XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[62]), .B (x[62]));
XOR2_X1 i_0_158 (.Z (u[63]), .A (z[62]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[50]), .A (z[50]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[49]), .B (x[62]));
XNOR2_X1 i_0_155 (.ZN (u[49]), .A (y[49]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_153 (.ZN (u[48]), .A (y[48]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_151 (.ZN (u[47]), .A (y[47]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_149 (.ZN (u[46]), .A (y[46]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_147 (.ZN (u[45]), .A (y[45]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_145 (.ZN (u[44]), .A (y[44]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_143 (.ZN (u[43]), .A (y[43]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_141 (.ZN (u[42]), .A (y[42]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_139 (.ZN (u[41]), .A (y[41]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_137 (.ZN (u[40]), .A (y[40]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_135 (.ZN (u[39]), .A (y[39]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_133 (.ZN (u[38]), .A (y[38]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_131 (.ZN (u[37]), .A (y[37]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_129 (.ZN (u[36]), .A (y[36]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_127 (.ZN (u[35]), .A (y[35]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_125 (.ZN (u[34]), .A (y[34]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_123 (.ZN (u[33]), .A (y[33]), .B (n_0_76));
XNOR2_X1 i_0_122 (.ZN (n_0_75), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_121 (.ZN (u[32]), .A (y[32]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_119 (.ZN (u[31]), .A (y[31]), .B (n_0_74));
XNOR2_X1 i_0_118 (.ZN (n_0_73), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_117 (.ZN (u[30]), .A (y[30]), .B (n_0_73));
XNOR2_X1 i_0_116 (.ZN (n_0_72), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_115 (.ZN (u[29]), .A (y[29]), .B (n_0_72));
XNOR2_X1 i_0_114 (.ZN (n_0_71), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_113 (.ZN (u[28]), .A (y[28]), .B (n_0_71));
XNOR2_X1 i_0_112 (.ZN (n_0_70), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_111 (.ZN (u[27]), .A (y[27]), .B (n_0_70));
XNOR2_X1 i_0_110 (.ZN (n_0_69), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_109 (.ZN (u[26]), .A (y[26]), .B (n_0_69));
XNOR2_X1 i_0_108 (.ZN (n_0_68), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_107 (.ZN (u[25]), .A (y[25]), .B (n_0_68));
XNOR2_X1 i_0_106 (.ZN (n_0_67), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_105 (.ZN (u[24]), .A (y[24]), .B (n_0_67));
XNOR2_X1 i_0_104 (.ZN (n_0_66), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_103 (.ZN (u[23]), .A (y[23]), .B (n_0_66));
XNOR2_X1 i_0_102 (.ZN (n_0_65), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_101 (.ZN (u[22]), .A (y[22]), .B (n_0_65));
XNOR2_X1 i_0_100 (.ZN (n_0_64), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_99 (.ZN (u[21]), .A (y[21]), .B (n_0_64));
XNOR2_X1 i_0_98 (.ZN (n_0_63), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_97 (.ZN (u[20]), .A (y[20]), .B (n_0_63));
XOR2_X1 i_0_96 (.Z (u[19]), .A (y[19]), .B (x[19]));
NAND2_X1 i_0_95 (.ZN (n_0_62), .A1 (y[62]), .A2 (x[62]));
OAI21_X1 i_0_94 (.ZN (n_0_61), .A (z[62]), .B1 (x[62]), .B2 (y[62]));
NAND2_X1 i_0_93 (.ZN (v[63]), .A1 (n_0_62), .A2 (n_0_61));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (z[50]), .B1 (x[62]), .B2 (y[62]));
NAND2_X1 i_0_91 (.ZN (v[51]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[49]), .A2 (x[62]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[49]), .B1 (z[49]), .B2 (x[62]));
NAND2_X1 i_0_88 (.ZN (v[50]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_85 (.ZN (v[49]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_82 (.ZN (v[48]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_79 (.ZN (v[47]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_76 (.ZN (v[46]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_73 (.ZN (v[45]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_70 (.ZN (v[44]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_67 (.ZN (v[43]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_64 (.ZN (v[42]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_61 (.ZN (v[41]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_58 (.ZN (v[40]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_55 (.ZN (v[39]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_52 (.ZN (v[38]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_49 (.ZN (v[37]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_46 (.ZN (v[36]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_43 (.ZN (v[35]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_40 (.ZN (v[34]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_37 (.ZN (v[33]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_34 (.ZN (v[32]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_31 (.ZN (v[31]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_28 (.ZN (v[30]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_25 (.ZN (v[29]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_22 (.ZN (v[28]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_19 (.ZN (v[27]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_16 (.ZN (v[26]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_13 (.ZN (v[25]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_10 (.ZN (v[24]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_7 (.ZN (v[23]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_4 (.ZN (v[22]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_1 (.ZN (v[21]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[20]), .A1 (y[19]), .A2 (x[19]));

endmodule //CSA__4_14

module CSA__4_11 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;


INV_X1 i_0_223 (.ZN (n_0_124), .A (x[62]));
INV_X1 i_0_222 (.ZN (n_0_123), .A (x[61]));
INV_X1 i_0_221 (.ZN (n_0_122), .A (x[60]));
INV_X1 i_0_220 (.ZN (n_0_121), .A (x[59]));
INV_X1 i_0_219 (.ZN (n_0_120), .A (x[58]));
INV_X1 i_0_218 (.ZN (n_0_119), .A (x[57]));
INV_X1 i_0_217 (.ZN (n_0_118), .A (x[56]));
INV_X1 i_0_216 (.ZN (n_0_117), .A (x[55]));
XOR2_X2 i_0_215 (.Z (n_0_116), .A (y[63]), .B (z[63]));
XOR2_X1 i_0_214 (.Z (u[63]), .A (x[63]), .B (n_0_116));
XNOR2_X1 i_0_213 (.ZN (u[62]), .A (n_0_124), .B (n_0_116));
XNOR2_X1 i_0_212 (.ZN (u[61]), .A (n_0_123), .B (n_0_116));
XNOR2_X1 i_0_211 (.ZN (u[60]), .A (n_0_122), .B (n_0_116));
XNOR2_X1 i_0_210 (.ZN (u[59]), .A (n_0_121), .B (n_0_116));
XNOR2_X1 i_0_209 (.ZN (u[58]), .A (n_0_120), .B (n_0_116));
XNOR2_X1 i_0_208 (.ZN (u[57]), .A (n_0_119), .B (n_0_116));
XNOR2_X1 i_0_207 (.ZN (u[56]), .A (n_0_118), .B (n_0_116));
XNOR2_X1 i_0_206 (.ZN (u[55]), .A (n_0_117), .B (n_0_116));
XNOR2_X1 i_0_205 (.ZN (n_0_115), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_204 (.ZN (u[54]), .A (y[63]), .B (n_0_115));
XNOR2_X1 i_0_203 (.ZN (n_0_114), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_202 (.ZN (u[53]), .A (y[53]), .B (n_0_114));
XNOR2_X1 i_0_201 (.ZN (n_0_113), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_200 (.ZN (u[52]), .A (y[52]), .B (n_0_113));
XNOR2_X1 i_0_199 (.ZN (n_0_112), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_198 (.ZN (u[51]), .A (y[51]), .B (n_0_112));
XNOR2_X1 i_0_197 (.ZN (n_0_111), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_196 (.ZN (u[50]), .A (y[50]), .B (n_0_111));
XNOR2_X1 i_0_195 (.ZN (n_0_110), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_194 (.ZN (u[49]), .A (y[49]), .B (n_0_110));
XNOR2_X1 i_0_193 (.ZN (n_0_109), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_192 (.ZN (u[48]), .A (y[48]), .B (n_0_109));
XNOR2_X1 i_0_191 (.ZN (n_0_108), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_190 (.ZN (u[47]), .A (y[47]), .B (n_0_108));
XNOR2_X1 i_0_189 (.ZN (n_0_107), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_188 (.ZN (u[46]), .A (y[46]), .B (n_0_107));
XNOR2_X1 i_0_187 (.ZN (n_0_106), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_186 (.ZN (u[45]), .A (y[45]), .B (n_0_106));
XNOR2_X1 i_0_185 (.ZN (n_0_105), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_184 (.ZN (u[44]), .A (y[44]), .B (n_0_105));
XNOR2_X1 i_0_183 (.ZN (n_0_104), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_182 (.ZN (u[43]), .A (y[43]), .B (n_0_104));
XNOR2_X1 i_0_181 (.ZN (n_0_103), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_180 (.ZN (u[42]), .A (y[42]), .B (n_0_103));
XNOR2_X1 i_0_179 (.ZN (n_0_102), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_178 (.ZN (u[41]), .A (y[41]), .B (n_0_102));
XNOR2_X1 i_0_177 (.ZN (n_0_101), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_176 (.ZN (u[40]), .A (y[40]), .B (n_0_101));
XNOR2_X1 i_0_175 (.ZN (n_0_100), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_174 (.ZN (u[39]), .A (y[39]), .B (n_0_100));
XNOR2_X1 i_0_173 (.ZN (n_0_99), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_172 (.ZN (u[38]), .A (y[38]), .B (n_0_99));
XNOR2_X1 i_0_171 (.ZN (n_0_98), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_170 (.ZN (u[37]), .A (y[37]), .B (n_0_98));
XNOR2_X1 i_0_169 (.ZN (n_0_97), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_168 (.ZN (u[36]), .A (y[36]), .B (n_0_97));
XNOR2_X1 i_0_167 (.ZN (n_0_96), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_166 (.ZN (u[35]), .A (y[35]), .B (n_0_96));
XNOR2_X1 i_0_165 (.ZN (n_0_95), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_164 (.ZN (u[34]), .A (y[34]), .B (n_0_95));
XNOR2_X1 i_0_163 (.ZN (n_0_94), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_162 (.ZN (u[33]), .A (y[33]), .B (n_0_94));
XNOR2_X1 i_0_161 (.ZN (n_0_93), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_160 (.ZN (u[32]), .A (y[32]), .B (n_0_93));
XNOR2_X1 i_0_159 (.ZN (n_0_92), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_158 (.ZN (u[31]), .A (y[31]), .B (n_0_92));
XNOR2_X1 i_0_157 (.ZN (n_0_91), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_156 (.ZN (u[30]), .A (y[30]), .B (n_0_91));
XNOR2_X1 i_0_155 (.ZN (n_0_90), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_154 (.ZN (u[29]), .A (y[29]), .B (n_0_90));
XNOR2_X1 i_0_153 (.ZN (n_0_89), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_152 (.ZN (u[28]), .A (y[28]), .B (n_0_89));
XNOR2_X1 i_0_151 (.ZN (n_0_88), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_150 (.ZN (u[27]), .A (y[27]), .B (n_0_88));
XNOR2_X1 i_0_149 (.ZN (n_0_87), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_148 (.ZN (u[26]), .A (y[26]), .B (n_0_87));
XNOR2_X1 i_0_147 (.ZN (n_0_86), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_146 (.ZN (u[25]), .A (y[25]), .B (n_0_86));
XNOR2_X1 i_0_145 (.ZN (n_0_85), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_144 (.ZN (u[24]), .A (y[24]), .B (n_0_85));
XNOR2_X1 i_0_143 (.ZN (n_0_84), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_142 (.ZN (u[23]), .A (y[23]), .B (n_0_84));
XNOR2_X1 i_0_141 (.ZN (n_0_83), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_140 (.ZN (u[22]), .A (y[22]), .B (n_0_83));
XNOR2_X1 i_0_139 (.ZN (n_0_82), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_138 (.ZN (u[21]), .A (y[21]), .B (n_0_82));
XNOR2_X1 i_0_137 (.ZN (n_0_81), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_136 (.ZN (u[20]), .A (y[20]), .B (n_0_81));
XNOR2_X1 i_0_135 (.ZN (n_0_80), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_134 (.ZN (u[19]), .A (y[19]), .B (n_0_80));
XNOR2_X1 i_0_133 (.ZN (n_0_79), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_132 (.ZN (u[18]), .A (y[18]), .B (n_0_79));
XNOR2_X1 i_0_131 (.ZN (n_0_78), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_130 (.ZN (u[17]), .A (y[17]), .B (n_0_78));
XOR2_X1 i_0_129 (.Z (u[16]), .A (y[16]), .B (x[16]));
XOR2_X1 i_0_128 (.Z (u[15]), .A (y[15]), .B (x[15]));
XOR2_X1 i_0_127 (.Z (u[14]), .A (y[14]), .B (x[14]));
NAND2_X1 i_0_126 (.ZN (n_0_77), .A1 (y[63]), .A2 (z[63]));
NOR2_X1 i_0_125 (.ZN (n_0_76), .A1 (y[63]), .A2 (z[63]));
OAI21_X1 i_0_124 (.ZN (v[63]), .A (n_0_77), .B1 (n_0_76), .B2 (n_0_124));
OAI21_X1 i_0_123 (.ZN (v[62]), .A (n_0_77), .B1 (n_0_76), .B2 (n_0_123));
OAI21_X1 i_0_122 (.ZN (v[61]), .A (n_0_77), .B1 (n_0_76), .B2 (n_0_122));
OAI21_X1 i_0_121 (.ZN (v[60]), .A (n_0_77), .B1 (n_0_76), .B2 (n_0_121));
OAI21_X1 i_0_120 (.ZN (v[59]), .A (n_0_77), .B1 (n_0_76), .B2 (n_0_120));
OAI21_X1 i_0_119 (.ZN (v[58]), .A (n_0_77), .B1 (n_0_76), .B2 (n_0_119));
OAI21_X1 i_0_118 (.ZN (v[57]), .A (n_0_77), .B1 (n_0_76), .B2 (n_0_118));
OAI21_X1 i_0_117 (.ZN (v[56]), .A (n_0_77), .B1 (n_0_76), .B2 (n_0_117));
NAND2_X1 i_0_116 (.ZN (n_0_75), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_115 (.ZN (n_0_74), .A (y[63]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_114 (.ZN (v[55]), .A1 (n_0_75), .A2 (n_0_74));
NAND2_X1 i_0_113 (.ZN (n_0_73), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_112 (.ZN (n_0_72), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_111 (.ZN (v[54]), .A1 (n_0_73), .A2 (n_0_72));
NAND2_X1 i_0_110 (.ZN (n_0_71), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_109 (.ZN (n_0_70), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_108 (.ZN (v[53]), .A1 (n_0_71), .A2 (n_0_70));
NAND2_X1 i_0_107 (.ZN (n_0_69), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_106 (.ZN (n_0_68), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_105 (.ZN (v[52]), .A1 (n_0_69), .A2 (n_0_68));
NAND2_X1 i_0_104 (.ZN (n_0_67), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_103 (.ZN (n_0_66), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_102 (.ZN (v[51]), .A1 (n_0_67), .A2 (n_0_66));
NAND2_X1 i_0_101 (.ZN (n_0_65), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_100 (.ZN (n_0_64), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_99 (.ZN (v[50]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_98 (.ZN (n_0_63), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_97 (.ZN (n_0_62), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_96 (.ZN (v[49]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_95 (.ZN (n_0_61), .A1 (y[47]), .A2 (x[47]));
OAI21_X1 i_0_94 (.ZN (n_0_60), .A (z[47]), .B1 (x[47]), .B2 (y[47]));
NAND2_X1 i_0_93 (.ZN (v[48]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_92 (.ZN (n_0_59), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_91 (.ZN (n_0_58), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_90 (.ZN (v[47]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_89 (.ZN (n_0_57), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_88 (.ZN (n_0_56), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_87 (.ZN (v[46]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_86 (.ZN (n_0_55), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_85 (.ZN (n_0_54), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_84 (.ZN (v[45]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_83 (.ZN (n_0_53), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_82 (.ZN (n_0_52), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_81 (.ZN (v[44]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_80 (.ZN (n_0_51), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_79 (.ZN (n_0_50), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_78 (.ZN (v[43]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_77 (.ZN (n_0_49), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_76 (.ZN (n_0_48), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_75 (.ZN (v[42]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_74 (.ZN (n_0_47), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_73 (.ZN (n_0_46), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_72 (.ZN (v[41]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_71 (.ZN (n_0_45), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_70 (.ZN (n_0_44), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_69 (.ZN (v[40]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_68 (.ZN (n_0_43), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_67 (.ZN (n_0_42), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_66 (.ZN (v[39]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_65 (.ZN (n_0_41), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_64 (.ZN (n_0_40), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_63 (.ZN (v[38]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_62 (.ZN (n_0_39), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_61 (.ZN (n_0_38), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_60 (.ZN (v[37]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_59 (.ZN (n_0_37), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_58 (.ZN (n_0_36), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_57 (.ZN (v[36]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_56 (.ZN (n_0_35), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_55 (.ZN (n_0_34), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_54 (.ZN (v[35]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_53 (.ZN (n_0_33), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_52 (.ZN (n_0_32), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_51 (.ZN (v[34]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_50 (.ZN (n_0_31), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_49 (.ZN (n_0_30), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_48 (.ZN (v[33]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_47 (.ZN (n_0_29), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_46 (.ZN (n_0_28), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_45 (.ZN (v[32]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_44 (.ZN (n_0_27), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_43 (.ZN (n_0_26), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_42 (.ZN (v[31]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_41 (.ZN (n_0_25), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_40 (.ZN (n_0_24), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_39 (.ZN (v[30]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_38 (.ZN (n_0_23), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_37 (.ZN (n_0_22), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_36 (.ZN (v[29]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_35 (.ZN (n_0_21), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_34 (.ZN (n_0_20), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_33 (.ZN (v[28]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_32 (.ZN (n_0_19), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_31 (.ZN (n_0_18), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_30 (.ZN (v[27]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_29 (.ZN (n_0_17), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_28 (.ZN (n_0_16), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_27 (.ZN (v[26]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_26 (.ZN (n_0_15), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_25 (.ZN (n_0_14), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_24 (.ZN (v[25]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_23 (.ZN (n_0_13), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_22 (.ZN (n_0_12), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_21 (.ZN (v[24]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_20 (.ZN (n_0_11), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_19 (.ZN (n_0_10), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_18 (.ZN (v[23]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_17 (.ZN (n_0_9), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_16 (.ZN (n_0_8), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_15 (.ZN (v[22]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_14 (.ZN (n_0_7), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_13 (.ZN (n_0_6), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_12 (.ZN (v[21]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_11 (.ZN (n_0_5), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_10 (.ZN (n_0_4), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_9 (.ZN (v[20]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_8 (.ZN (n_0_3), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_7 (.ZN (n_0_2), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_6 (.ZN (v[19]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_5 (.ZN (n_0_1), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_4 (.ZN (n_0_0), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_3 (.ZN (v[18]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_2 (.ZN (v[17]), .A1 (y[16]), .A2 (x[16]));
AND2_X1 i_0_1 (.ZN (v[16]), .A1 (y[15]), .A2 (x[15]));
AND2_X1 i_0_0 (.ZN (v[15]), .A1 (y[14]), .A2 (x[14]));

endmodule //CSA__4_11

module CSA__4_8 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;


INV_X1 i_0_181 (.ZN (n_0_103), .A (z[63]));
INV_X1 i_0_180 (.ZN (n_0_102), .A (z[53]));
INV_X1 i_0_179 (.ZN (n_0_101), .A (z[52]));
INV_X1 i_0_178 (.ZN (n_0_100), .A (z[51]));
INV_X1 i_0_177 (.ZN (n_0_99), .A (z[50]));
XOR2_X1 i_0_176 (.Z (n_0_98), .A (y[63]), .B (x[63]));
XNOR2_X1 i_0_175 (.ZN (u[63]), .A (n_0_103), .B (n_0_98));
XNOR2_X1 i_0_174 (.ZN (u[53]), .A (n_0_102), .B (n_0_98));
XNOR2_X1 i_0_173 (.ZN (u[52]), .A (n_0_101), .B (n_0_98));
XNOR2_X1 i_0_172 (.ZN (u[51]), .A (n_0_100), .B (n_0_98));
XNOR2_X1 i_0_171 (.ZN (u[50]), .A (n_0_99), .B (n_0_98));
XNOR2_X1 i_0_170 (.ZN (n_0_97), .A (z[49]), .B (x[63]));
XNOR2_X1 i_0_169 (.ZN (u[49]), .A (y[49]), .B (n_0_97));
XNOR2_X1 i_0_168 (.ZN (n_0_96), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_167 (.ZN (u[48]), .A (y[48]), .B (n_0_96));
XNOR2_X1 i_0_166 (.ZN (n_0_95), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_165 (.ZN (u[47]), .A (y[47]), .B (n_0_95));
XNOR2_X1 i_0_164 (.ZN (n_0_94), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_163 (.ZN (u[46]), .A (y[46]), .B (n_0_94));
XNOR2_X1 i_0_162 (.ZN (n_0_93), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_161 (.ZN (u[45]), .A (y[45]), .B (n_0_93));
XNOR2_X1 i_0_160 (.ZN (n_0_92), .A (z[44]), .B (x[44]));
XNOR2_X2 i_0_159 (.ZN (u[44]), .A (y[44]), .B (n_0_92));
XNOR2_X1 i_0_158 (.ZN (n_0_91), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_157 (.ZN (u[43]), .A (y[43]), .B (n_0_91));
XNOR2_X1 i_0_156 (.ZN (n_0_90), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_155 (.ZN (u[42]), .A (y[42]), .B (n_0_90));
XNOR2_X1 i_0_154 (.ZN (n_0_89), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_153 (.ZN (u[41]), .A (y[41]), .B (n_0_89));
XNOR2_X1 i_0_152 (.ZN (n_0_88), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_151 (.ZN (u[40]), .A (y[40]), .B (n_0_88));
XNOR2_X1 i_0_150 (.ZN (n_0_87), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_149 (.ZN (u[39]), .A (y[39]), .B (n_0_87));
XNOR2_X1 i_0_148 (.ZN (n_0_86), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_147 (.ZN (u[38]), .A (y[38]), .B (n_0_86));
XNOR2_X1 i_0_146 (.ZN (n_0_85), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_145 (.ZN (u[37]), .A (y[37]), .B (n_0_85));
XNOR2_X1 i_0_144 (.ZN (n_0_84), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_143 (.ZN (u[36]), .A (y[36]), .B (n_0_84));
XNOR2_X1 i_0_142 (.ZN (n_0_83), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_141 (.ZN (u[35]), .A (y[35]), .B (n_0_83));
XNOR2_X1 i_0_140 (.ZN (n_0_82), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_139 (.ZN (u[34]), .A (y[34]), .B (n_0_82));
XNOR2_X1 i_0_138 (.ZN (n_0_81), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_137 (.ZN (u[33]), .A (y[33]), .B (n_0_81));
XNOR2_X1 i_0_136 (.ZN (n_0_80), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_135 (.ZN (u[32]), .A (y[32]), .B (n_0_80));
XNOR2_X1 i_0_134 (.ZN (n_0_79), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_133 (.ZN (u[31]), .A (y[31]), .B (n_0_79));
XNOR2_X1 i_0_132 (.ZN (n_0_78), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_131 (.ZN (u[30]), .A (y[30]), .B (n_0_78));
XNOR2_X1 i_0_130 (.ZN (n_0_77), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_129 (.ZN (u[29]), .A (y[29]), .B (n_0_77));
XNOR2_X1 i_0_128 (.ZN (n_0_76), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_127 (.ZN (u[28]), .A (y[28]), .B (n_0_76));
XNOR2_X1 i_0_126 (.ZN (n_0_75), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_125 (.ZN (u[27]), .A (y[27]), .B (n_0_75));
XNOR2_X1 i_0_124 (.ZN (n_0_74), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_123 (.ZN (u[26]), .A (y[26]), .B (n_0_74));
XNOR2_X1 i_0_122 (.ZN (n_0_73), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_121 (.ZN (u[25]), .A (y[25]), .B (n_0_73));
XNOR2_X1 i_0_120 (.ZN (n_0_72), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_119 (.ZN (u[24]), .A (y[24]), .B (n_0_72));
XNOR2_X1 i_0_118 (.ZN (n_0_71), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_117 (.ZN (u[23]), .A (y[23]), .B (n_0_71));
XNOR2_X1 i_0_116 (.ZN (n_0_70), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_115 (.ZN (u[22]), .A (y[22]), .B (n_0_70));
XNOR2_X1 i_0_114 (.ZN (n_0_69), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_113 (.ZN (u[21]), .A (y[21]), .B (n_0_69));
XNOR2_X1 i_0_112 (.ZN (n_0_68), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_111 (.ZN (u[20]), .A (y[20]), .B (n_0_68));
XNOR2_X1 i_0_110 (.ZN (n_0_67), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_109 (.ZN (u[19]), .A (y[19]), .B (n_0_67));
XNOR2_X1 i_0_108 (.ZN (n_0_66), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_107 (.ZN (u[18]), .A (y[18]), .B (n_0_66));
XOR2_X1 i_0_106 (.Z (u[17]), .A (y[17]), .B (x[17]));
XOR2_X1 i_0_105 (.Z (u[16]), .A (y[16]), .B (x[16]));
NOR2_X1 i_0_104 (.ZN (n_0_65), .A1 (y[63]), .A2 (x[63]));
NAND2_X1 i_0_103 (.ZN (n_0_64), .A1 (y[63]), .A2 (x[63]));
AOI21_X1 i_0_102 (.ZN (v[63]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_103));
AOI21_X1 i_0_101 (.ZN (v[54]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_102));
AOI21_X1 i_0_100 (.ZN (v[53]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_101));
AOI21_X1 i_0_99 (.ZN (v[52]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_100));
AOI21_X1 i_0_98 (.ZN (v[51]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_99));
NAND2_X1 i_0_97 (.ZN (n_0_63), .A1 (z[49]), .A2 (x[63]));
OAI21_X1 i_0_96 (.ZN (n_0_62), .A (y[49]), .B1 (z[49]), .B2 (x[63]));
NAND2_X1 i_0_95 (.ZN (v[50]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_94 (.ZN (n_0_61), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_93 (.ZN (n_0_60), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_92 (.ZN (v[49]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_91 (.ZN (n_0_59), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_90 (.ZN (n_0_58), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_89 (.ZN (v[48]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_88 (.ZN (n_0_57), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_87 (.ZN (n_0_56), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_86 (.ZN (v[47]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_85 (.ZN (n_0_55), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_84 (.ZN (n_0_54), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_83 (.ZN (v[46]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_82 (.ZN (n_0_53), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_81 (.ZN (n_0_52), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_80 (.ZN (v[45]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_79 (.ZN (n_0_51), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_78 (.ZN (n_0_50), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_77 (.ZN (v[44]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_76 (.ZN (n_0_49), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_75 (.ZN (n_0_48), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_74 (.ZN (v[43]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_73 (.ZN (n_0_47), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_72 (.ZN (n_0_46), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_71 (.ZN (v[42]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_70 (.ZN (n_0_45), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_69 (.ZN (n_0_44), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_68 (.ZN (v[41]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_67 (.ZN (n_0_43), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_66 (.ZN (n_0_42), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_65 (.ZN (v[40]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_64 (.ZN (n_0_41), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_63 (.ZN (n_0_40), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_62 (.ZN (v[39]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_61 (.ZN (n_0_39), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_60 (.ZN (n_0_38), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_59 (.ZN (v[38]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_58 (.ZN (n_0_37), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_57 (.ZN (n_0_36), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_56 (.ZN (v[37]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_55 (.ZN (n_0_35), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_54 (.ZN (n_0_34), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_53 (.ZN (v[36]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_52 (.ZN (n_0_33), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_51 (.ZN (n_0_32), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_50 (.ZN (v[35]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_49 (.ZN (n_0_31), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_48 (.ZN (n_0_30), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_47 (.ZN (v[34]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_46 (.ZN (n_0_29), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_45 (.ZN (n_0_28), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_44 (.ZN (v[33]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_43 (.ZN (n_0_27), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_42 (.ZN (n_0_26), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_41 (.ZN (v[32]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_40 (.ZN (n_0_25), .A1 (y[30]), .A2 (z[30]));
OAI21_X1 i_0_39 (.ZN (n_0_24), .A (x[30]), .B1 (z[30]), .B2 (y[30]));
NAND2_X1 i_0_38 (.ZN (v[31]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_37 (.ZN (n_0_23), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_36 (.ZN (n_0_22), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_35 (.ZN (v[30]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_34 (.ZN (n_0_21), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_33 (.ZN (n_0_20), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_32 (.ZN (v[29]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_31 (.ZN (n_0_19), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_30 (.ZN (n_0_18), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_29 (.ZN (v[28]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_28 (.ZN (n_0_17), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_27 (.ZN (n_0_16), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_26 (.ZN (v[27]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_25 (.ZN (n_0_15), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_24 (.ZN (n_0_14), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_23 (.ZN (v[26]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_22 (.ZN (n_0_13), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_21 (.ZN (n_0_12), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_20 (.ZN (v[25]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_19 (.ZN (n_0_11), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_18 (.ZN (n_0_10), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_17 (.ZN (v[24]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_16 (.ZN (n_0_9), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_15 (.ZN (n_0_8), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_14 (.ZN (v[23]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_13 (.ZN (n_0_7), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_12 (.ZN (n_0_6), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_11 (.ZN (v[22]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_10 (.ZN (n_0_5), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_9 (.ZN (n_0_4), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_8 (.ZN (v[21]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_7 (.ZN (n_0_3), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_6 (.ZN (n_0_2), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_5 (.ZN (v[20]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_4 (.ZN (n_0_1), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_3 (.ZN (n_0_0), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_2 (.ZN (v[19]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_1 (.ZN (v[18]), .A1 (y[17]), .A2 (x[17]));
AND2_X1 i_0_0 (.ZN (v[17]), .A1 (y[16]), .A2 (x[16]));

endmodule //CSA__4_8

module CSA__4_5 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;


INV_X1 i_0_168 (.ZN (n_0_98), .A (z[63]));
INV_X1 i_0_167 (.ZN (n_0_97), .A (z[53]));
INV_X1 i_0_166 (.ZN (n_0_96), .A (z[52]));
XOR2_X1 i_0_165 (.Z (n_0_95), .A (y[63]), .B (x[63]));
XNOR2_X1 i_0_164 (.ZN (u[63]), .A (n_0_98), .B (n_0_95));
XNOR2_X1 i_0_163 (.ZN (u[53]), .A (n_0_97), .B (n_0_95));
XNOR2_X1 i_0_162 (.ZN (u[52]), .A (n_0_96), .B (n_0_95));
XNOR2_X1 i_0_161 (.ZN (n_0_94), .A (z[51]), .B (x[63]));
XNOR2_X1 i_0_160 (.ZN (u[51]), .A (y[51]), .B (n_0_94));
XNOR2_X1 i_0_159 (.ZN (n_0_93), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_158 (.ZN (u[50]), .A (y[50]), .B (n_0_93));
XNOR2_X1 i_0_157 (.ZN (n_0_92), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_156 (.ZN (u[49]), .A (y[49]), .B (n_0_92));
XNOR2_X1 i_0_155 (.ZN (n_0_91), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_154 (.ZN (u[48]), .A (y[48]), .B (n_0_91));
XNOR2_X1 i_0_153 (.ZN (n_0_90), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_152 (.ZN (u[47]), .A (y[47]), .B (n_0_90));
XNOR2_X1 i_0_151 (.ZN (n_0_89), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_150 (.ZN (u[46]), .A (y[46]), .B (n_0_89));
XNOR2_X1 i_0_149 (.ZN (n_0_88), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_148 (.ZN (u[45]), .A (y[45]), .B (n_0_88));
XNOR2_X1 i_0_147 (.ZN (n_0_87), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_146 (.ZN (u[44]), .A (y[44]), .B (n_0_87));
XNOR2_X1 i_0_145 (.ZN (n_0_86), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_144 (.ZN (u[43]), .A (y[43]), .B (n_0_86));
XNOR2_X1 i_0_143 (.ZN (n_0_85), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_142 (.ZN (u[42]), .A (y[42]), .B (n_0_85));
XNOR2_X1 i_0_141 (.ZN (n_0_84), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_140 (.ZN (u[41]), .A (y[41]), .B (n_0_84));
XNOR2_X1 i_0_139 (.ZN (n_0_83), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_138 (.ZN (u[40]), .A (y[40]), .B (n_0_83));
XNOR2_X1 i_0_137 (.ZN (n_0_82), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_136 (.ZN (u[39]), .A (y[39]), .B (n_0_82));
XNOR2_X1 i_0_135 (.ZN (n_0_81), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_134 (.ZN (u[38]), .A (y[38]), .B (n_0_81));
XNOR2_X1 i_0_133 (.ZN (n_0_80), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_132 (.ZN (u[37]), .A (y[37]), .B (n_0_80));
XNOR2_X1 i_0_131 (.ZN (n_0_79), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_130 (.ZN (u[36]), .A (y[36]), .B (n_0_79));
XNOR2_X1 i_0_129 (.ZN (n_0_78), .A (z[35]), .B (x[35]));
XNOR2_X2 i_0_128 (.ZN (u[35]), .A (y[35]), .B (n_0_78));
XNOR2_X1 i_0_127 (.ZN (n_0_77), .A (z[34]), .B (x[34]));
XNOR2_X2 i_0_126 (.ZN (u[34]), .A (y[34]), .B (n_0_77));
XNOR2_X1 i_0_125 (.ZN (n_0_76), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_124 (.ZN (u[33]), .A (y[33]), .B (n_0_76));
XNOR2_X1 i_0_123 (.ZN (n_0_75), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_122 (.ZN (u[32]), .A (y[32]), .B (n_0_75));
XNOR2_X1 i_0_121 (.ZN (n_0_74), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_120 (.ZN (u[31]), .A (y[31]), .B (n_0_74));
XNOR2_X1 i_0_119 (.ZN (n_0_73), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_118 (.ZN (u[30]), .A (y[30]), .B (n_0_73));
XNOR2_X1 i_0_117 (.ZN (n_0_72), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_116 (.ZN (u[29]), .A (y[29]), .B (n_0_72));
XNOR2_X1 i_0_115 (.ZN (n_0_71), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_114 (.ZN (u[28]), .A (y[28]), .B (n_0_71));
XNOR2_X1 i_0_113 (.ZN (n_0_70), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_112 (.ZN (u[27]), .A (y[27]), .B (n_0_70));
XNOR2_X1 i_0_111 (.ZN (n_0_69), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_110 (.ZN (u[26]), .A (y[26]), .B (n_0_69));
XNOR2_X1 i_0_109 (.ZN (n_0_68), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_108 (.ZN (u[25]), .A (y[25]), .B (n_0_68));
XNOR2_X1 i_0_107 (.ZN (n_0_67), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_106 (.ZN (u[24]), .A (y[24]), .B (n_0_67));
XNOR2_X1 i_0_105 (.ZN (n_0_66), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_104 (.ZN (u[23]), .A (y[23]), .B (n_0_66));
XNOR2_X1 i_0_103 (.ZN (n_0_65), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_102 (.ZN (u[22]), .A (y[22]), .B (n_0_65));
XNOR2_X1 i_0_101 (.ZN (n_0_64), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_100 (.ZN (u[21]), .A (y[21]), .B (n_0_64));
XOR2_X1 i_0_99 (.Z (u[20]), .A (y[20]), .B (x[20]));
NOR2_X1 i_0_98 (.ZN (n_0_63), .A1 (y[63]), .A2 (x[63]));
NAND2_X1 i_0_97 (.ZN (n_0_62), .A1 (y[63]), .A2 (x[63]));
AOI21_X2 i_0_96 (.ZN (v[63]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_98));
AOI21_X1 i_0_95 (.ZN (v[54]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_97));
AOI21_X1 i_0_94 (.ZN (v[53]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_96));
NAND2_X1 i_0_93 (.ZN (n_0_61), .A1 (z[51]), .A2 (x[63]));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (y[51]), .B1 (z[51]), .B2 (x[63]));
NAND2_X1 i_0_91 (.ZN (v[52]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_88 (.ZN (v[51]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_85 (.ZN (v[50]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_82 (.ZN (v[49]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_79 (.ZN (v[48]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_76 (.ZN (v[47]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_73 (.ZN (v[46]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_70 (.ZN (v[45]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_67 (.ZN (v[44]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_64 (.ZN (v[43]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_61 (.ZN (v[42]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_58 (.ZN (v[41]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_55 (.ZN (v[40]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_52 (.ZN (v[39]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_49 (.ZN (v[38]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_46 (.ZN (v[37]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_43 (.ZN (v[36]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_40 (.ZN (v[35]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_37 (.ZN (v[34]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_34 (.ZN (v[33]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_31 (.ZN (v[32]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_28 (.ZN (v[31]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_25 (.ZN (v[30]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_22 (.ZN (v[29]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_19 (.ZN (v[28]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_16 (.ZN (v[27]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_13 (.ZN (v[26]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_10 (.ZN (v[25]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_7 (.ZN (v[24]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_4 (.ZN (v[23]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_1 (.ZN (v[22]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[21]), .A1 (y[20]), .A2 (x[20]));

endmodule //CSA__4_5

module CSA__4_2 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;


XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[63]), .B (x[63]));
XOR2_X1 i_0_158 (.Z (u[63]), .A (z[63]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[53]), .A (z[53]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[52]), .B (x[63]));
XNOR2_X1 i_0_155 (.ZN (u[52]), .A (y[52]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_153 (.ZN (u[51]), .A (y[51]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_151 (.ZN (u[50]), .A (y[50]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_149 (.ZN (u[49]), .A (y[49]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_147 (.ZN (u[48]), .A (y[48]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_145 (.ZN (u[47]), .A (y[47]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_143 (.ZN (u[46]), .A (y[46]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_141 (.ZN (u[45]), .A (y[45]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_139 (.ZN (u[44]), .A (y[44]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_137 (.ZN (u[43]), .A (y[43]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_135 (.ZN (u[42]), .A (y[42]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_133 (.ZN (u[41]), .A (y[41]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_131 (.ZN (u[40]), .A (y[40]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_129 (.ZN (u[39]), .A (y[39]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_127 (.ZN (u[38]), .A (y[38]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_125 (.ZN (u[37]), .A (y[37]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_123 (.ZN (u[36]), .A (y[36]), .B (n_0_76));
XNOR2_X1 i_0_122 (.ZN (n_0_75), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_121 (.ZN (u[35]), .A (y[35]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_119 (.ZN (u[34]), .A (y[34]), .B (n_0_74));
XNOR2_X1 i_0_118 (.ZN (n_0_73), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_117 (.ZN (u[33]), .A (y[33]), .B (n_0_73));
XNOR2_X1 i_0_116 (.ZN (n_0_72), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_115 (.ZN (u[32]), .A (y[32]), .B (n_0_72));
XNOR2_X1 i_0_114 (.ZN (n_0_71), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_113 (.ZN (u[31]), .A (y[31]), .B (n_0_71));
XNOR2_X1 i_0_112 (.ZN (n_0_70), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_111 (.ZN (u[30]), .A (y[30]), .B (n_0_70));
XNOR2_X1 i_0_110 (.ZN (n_0_69), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_109 (.ZN (u[29]), .A (y[29]), .B (n_0_69));
XNOR2_X1 i_0_108 (.ZN (n_0_68), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_107 (.ZN (u[28]), .A (y[28]), .B (n_0_68));
XNOR2_X1 i_0_106 (.ZN (n_0_67), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_105 (.ZN (u[27]), .A (y[27]), .B (n_0_67));
XNOR2_X1 i_0_104 (.ZN (n_0_66), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_103 (.ZN (u[26]), .A (y[26]), .B (n_0_66));
XNOR2_X1 i_0_102 (.ZN (n_0_65), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_101 (.ZN (u[25]), .A (y[25]), .B (n_0_65));
XNOR2_X1 i_0_100 (.ZN (n_0_64), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_99 (.ZN (u[24]), .A (y[24]), .B (n_0_64));
XNOR2_X1 i_0_98 (.ZN (n_0_63), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_97 (.ZN (u[23]), .A (y[23]), .B (n_0_63));
XOR2_X1 i_0_96 (.Z (u[22]), .A (y[22]), .B (x[22]));
NAND2_X1 i_0_95 (.ZN (n_0_62), .A1 (y[63]), .A2 (x[63]));
OAI21_X1 i_0_94 (.ZN (n_0_61), .A (z[63]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_93 (.ZN (v[63]), .A1 (n_0_62), .A2 (n_0_61));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (z[53]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_91 (.ZN (v[54]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[52]), .A2 (x[63]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[52]), .B1 (z[52]), .B2 (x[63]));
NAND2_X1 i_0_88 (.ZN (v[53]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_85 (.ZN (v[52]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_82 (.ZN (v[51]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_79 (.ZN (v[50]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_76 (.ZN (v[49]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_73 (.ZN (v[48]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_70 (.ZN (v[47]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_67 (.ZN (v[46]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_64 (.ZN (v[45]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_61 (.ZN (v[44]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_58 (.ZN (v[43]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_55 (.ZN (v[42]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_52 (.ZN (v[41]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_49 (.ZN (v[40]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_46 (.ZN (v[39]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_43 (.ZN (v[38]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_40 (.ZN (v[37]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_37 (.ZN (v[36]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_34 (.ZN (v[35]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_31 (.ZN (v[34]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_28 (.ZN (v[33]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_25 (.ZN (v[32]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_22 (.ZN (v[31]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_19 (.ZN (v[30]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_16 (.ZN (v[29]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_13 (.ZN (v[28]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_10 (.ZN (v[27]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_7 (.ZN (v[26]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_4 (.ZN (v[25]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_1 (.ZN (v[24]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[23]), .A1 (y[22]), .A2 (x[22]));

endmodule //CSA__4_2

module CSA__0_75 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire slo__mro_n7;


XNOR2_X1 i_0_276 (.ZN (n_0_159), .A (z[63]), .B (x[63]));
XNOR2_X1 i_0_275 (.ZN (u[63]), .A (y[63]), .B (n_0_159));
XNOR2_X1 i_0_274 (.ZN (n_0_158), .A (z[62]), .B (x[62]));
XNOR2_X1 i_0_273 (.ZN (u[62]), .A (y[62]), .B (n_0_158));
XNOR2_X1 i_0_272 (.ZN (n_0_157), .A (z[61]), .B (x[61]));
XNOR2_X1 i_0_271 (.ZN (u[61]), .A (y[61]), .B (n_0_157));
XNOR2_X1 i_0_270 (.ZN (n_0_156), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_269 (.ZN (u[60]), .A (y[60]), .B (n_0_156));
XNOR2_X1 i_0_268 (.ZN (n_0_155), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_267 (.ZN (u[59]), .A (y[59]), .B (n_0_155));
XNOR2_X1 i_0_266 (.ZN (n_0_154), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_265 (.ZN (u[58]), .A (y[58]), .B (n_0_154));
XNOR2_X1 i_0_264 (.ZN (n_0_153), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_263 (.ZN (u[57]), .A (y[57]), .B (n_0_153));
XNOR2_X1 i_0_262 (.ZN (n_0_152), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_261 (.ZN (u[56]), .A (y[56]), .B (n_0_152));
XNOR2_X1 i_0_260 (.ZN (n_0_151), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_259 (.ZN (u[55]), .A (y[55]), .B (n_0_151));
XNOR2_X1 i_0_258 (.ZN (n_0_150), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_257 (.ZN (u[54]), .A (y[54]), .B (n_0_150));
XNOR2_X1 i_0_256 (.ZN (n_0_149), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_255 (.ZN (u[53]), .A (y[53]), .B (n_0_149));
XNOR2_X1 i_0_254 (.ZN (n_0_148), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_253 (.ZN (u[52]), .A (y[52]), .B (n_0_148));
XNOR2_X1 i_0_252 (.ZN (n_0_147), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_251 (.ZN (u[51]), .A (y[51]), .B (n_0_147));
XNOR2_X1 i_0_250 (.ZN (n_0_146), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_249 (.ZN (u[50]), .A (y[50]), .B (n_0_146));
XNOR2_X1 i_0_248 (.ZN (n_0_145), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_247 (.ZN (u[49]), .A (y[49]), .B (n_0_145));
XNOR2_X1 i_0_246 (.ZN (n_0_144), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_245 (.ZN (u[48]), .A (y[48]), .B (n_0_144));
XNOR2_X1 i_0_244 (.ZN (n_0_143), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_243 (.ZN (u[47]), .A (y[47]), .B (n_0_143));
XNOR2_X1 i_0_242 (.ZN (n_0_142), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_241 (.ZN (u[46]), .A (y[46]), .B (n_0_142));
XNOR2_X1 i_0_240 (.ZN (n_0_141), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_239 (.ZN (u[45]), .A (y[45]), .B (n_0_141));
XNOR2_X1 i_0_238 (.ZN (n_0_140), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_237 (.ZN (u[44]), .A (y[44]), .B (n_0_140));
XNOR2_X1 i_0_236 (.ZN (n_0_139), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_235 (.ZN (u[43]), .A (y[43]), .B (n_0_139));
XNOR2_X1 i_0_234 (.ZN (n_0_138), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_233 (.ZN (u[42]), .A (y[42]), .B (n_0_138));
XNOR2_X1 i_0_232 (.ZN (n_0_137), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_231 (.ZN (u[41]), .A (y[41]), .B (n_0_137));
XNOR2_X1 i_0_230 (.ZN (n_0_136), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_229 (.ZN (u[40]), .A (y[40]), .B (n_0_136));
XNOR2_X1 i_0_228 (.ZN (n_0_135), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_227 (.ZN (u[39]), .A (y[39]), .B (n_0_135));
XNOR2_X1 i_0_226 (.ZN (n_0_134), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_225 (.ZN (u[38]), .A (y[38]), .B (n_0_134));
XNOR2_X1 i_0_224 (.ZN (n_0_133), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_223 (.ZN (u[37]), .A (y[37]), .B (n_0_133));
XNOR2_X1 i_0_222 (.ZN (n_0_132), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_221 (.ZN (u[36]), .A (y[36]), .B (n_0_132));
XNOR2_X1 i_0_220 (.ZN (n_0_131), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_219 (.ZN (u[35]), .A (y[35]), .B (n_0_131));
XNOR2_X1 i_0_218 (.ZN (n_0_130), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_217 (.ZN (u[34]), .A (y[34]), .B (n_0_130));
XNOR2_X1 i_0_216 (.ZN (n_0_129), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_215 (.ZN (u[33]), .A (y[33]), .B (n_0_129));
XNOR2_X1 i_0_214 (.ZN (n_0_128), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_213 (.ZN (u[32]), .A (y[32]), .B (n_0_128));
XNOR2_X1 i_0_212 (.ZN (n_0_127), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_211 (.ZN (u[31]), .A (y[31]), .B (n_0_127));
XNOR2_X1 i_0_210 (.ZN (n_0_126), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_209 (.ZN (u[30]), .A (y[30]), .B (n_0_126));
XNOR2_X1 i_0_208 (.ZN (n_0_125), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_207 (.ZN (u[29]), .A (y[29]), .B (n_0_125));
XNOR2_X1 i_0_206 (.ZN (n_0_124), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_205 (.ZN (u[28]), .A (y[28]), .B (n_0_124));
XNOR2_X1 i_0_204 (.ZN (n_0_123), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_203 (.ZN (u[27]), .A (y[27]), .B (n_0_123));
XNOR2_X1 i_0_202 (.ZN (n_0_122), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_201 (.ZN (u[26]), .A (y[26]), .B (n_0_122));
XNOR2_X1 i_0_200 (.ZN (n_0_121), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_199 (.ZN (u[25]), .A (y[25]), .B (n_0_121));
XNOR2_X1 i_0_198 (.ZN (n_0_120), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_197 (.ZN (u[24]), .A (y[24]), .B (n_0_120));
XNOR2_X1 i_0_196 (.ZN (n_0_119), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_195 (.ZN (u[23]), .A (y[23]), .B (n_0_119));
XNOR2_X1 i_0_194 (.ZN (n_0_118), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_193 (.ZN (u[22]), .A (y[22]), .B (n_0_118));
XNOR2_X1 i_0_192 (.ZN (n_0_117), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_191 (.ZN (u[21]), .A (y[21]), .B (n_0_117));
XNOR2_X1 i_0_190 (.ZN (n_0_116), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_189 (.ZN (u[20]), .A (y[20]), .B (n_0_116));
XNOR2_X1 i_0_188 (.ZN (n_0_115), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_187 (.ZN (u[19]), .A (y[19]), .B (n_0_115));
XNOR2_X1 i_0_186 (.ZN (n_0_114), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_185 (.ZN (u[18]), .A (y[18]), .B (n_0_114));
XNOR2_X1 i_0_184 (.ZN (n_0_113), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_183 (.ZN (u[17]), .A (y[17]), .B (n_0_113));
XNOR2_X2 i_0_182 (.ZN (n_0_112), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_181 (.ZN (u[16]), .A (y[16]), .B (n_0_112));
XNOR2_X2 i_0_180 (.ZN (n_0_111), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_179 (.ZN (u[15]), .A (n_0_111), .B (y[15]));
XNOR2_X2 i_0_178 (.ZN (n_0_110), .A (z[14]), .B (x[14]));
XNOR2_X2 i_0_177 (.ZN (u[14]), .A (y[14]), .B (n_0_110));
XNOR2_X2 i_0_174 (.ZN (n_0_108), .A (x[12]), .B (z[12]));
XNOR2_X2 i_0_173 (.ZN (u[12]), .A (n_0_108), .B (y[12]));
XNOR2_X2 i_0_172 (.ZN (n_0_107), .A (x[11]), .B (z[11]));
XNOR2_X2 i_0_171 (.ZN (u[11]), .A (n_0_107), .B (y[11]));
XNOR2_X2 i_0_170 (.ZN (n_0_106), .A (x[10]), .B (z[10]));
XNOR2_X2 i_0_169 (.ZN (u[10]), .A (n_0_106), .B (y[10]));
XOR2_X2 i_0_168 (.Z (u[9]), .A (y[9]), .B (x[9]));
XOR2_X2 i_0_167 (.Z (u[8]), .A (y[8]), .B (x[8]));
XOR2_X2 i_0_166 (.Z (u[7]), .A (y[7]), .B (x[7]));
XOR2_X1 i_0_165 (.Z (u[6]), .A (y[6]), .B (x[6]));
XOR2_X1 i_0_164 (.Z (u[5]), .A (y[5]), .B (x[5]));
NAND2_X1 i_0_163 (.ZN (n_0_105), .A1 (z[62]), .A2 (x[62]));
OAI21_X1 i_0_162 (.ZN (n_0_104), .A (y[62]), .B1 (z[62]), .B2 (x[62]));
NAND2_X1 i_0_161 (.ZN (v[63]), .A1 (n_0_105), .A2 (n_0_104));
NAND2_X1 i_0_160 (.ZN (n_0_103), .A1 (z[61]), .A2 (x[61]));
OAI21_X1 i_0_159 (.ZN (n_0_102), .A (y[61]), .B1 (z[61]), .B2 (x[61]));
NAND2_X1 i_0_158 (.ZN (v[62]), .A1 (n_0_103), .A2 (n_0_102));
NAND2_X1 i_0_157 (.ZN (n_0_101), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_156 (.ZN (n_0_100), .A (y[60]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_155 (.ZN (v[61]), .A1 (n_0_101), .A2 (n_0_100));
NAND2_X1 i_0_154 (.ZN (n_0_99), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_153 (.ZN (n_0_98), .A (y[59]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_152 (.ZN (v[60]), .A1 (n_0_99), .A2 (n_0_98));
NAND2_X1 i_0_151 (.ZN (n_0_97), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_150 (.ZN (n_0_96), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_149 (.ZN (v[59]), .A1 (n_0_97), .A2 (n_0_96));
NAND2_X1 i_0_148 (.ZN (n_0_95), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_147 (.ZN (n_0_94), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_146 (.ZN (v[58]), .A1 (n_0_95), .A2 (n_0_94));
NAND2_X1 i_0_145 (.ZN (n_0_93), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_144 (.ZN (n_0_92), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_143 (.ZN (v[57]), .A1 (n_0_93), .A2 (n_0_92));
NAND2_X1 i_0_142 (.ZN (n_0_91), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_141 (.ZN (n_0_90), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_140 (.ZN (v[56]), .A1 (n_0_91), .A2 (n_0_90));
NAND2_X1 i_0_139 (.ZN (n_0_89), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_138 (.ZN (n_0_88), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_137 (.ZN (v[55]), .A1 (n_0_89), .A2 (n_0_88));
NAND2_X1 i_0_136 (.ZN (n_0_87), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_135 (.ZN (n_0_86), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_134 (.ZN (v[54]), .A1 (n_0_87), .A2 (n_0_86));
NAND2_X1 i_0_133 (.ZN (n_0_85), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_132 (.ZN (n_0_84), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_131 (.ZN (v[53]), .A1 (n_0_85), .A2 (n_0_84));
NAND2_X1 i_0_130 (.ZN (n_0_83), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_129 (.ZN (n_0_82), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_128 (.ZN (v[52]), .A1 (n_0_83), .A2 (n_0_82));
NAND2_X1 i_0_127 (.ZN (n_0_81), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_126 (.ZN (n_0_80), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_125 (.ZN (v[51]), .A1 (n_0_81), .A2 (n_0_80));
NAND2_X1 i_0_124 (.ZN (n_0_79), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_123 (.ZN (n_0_78), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_122 (.ZN (v[50]), .A1 (n_0_79), .A2 (n_0_78));
NAND2_X1 i_0_121 (.ZN (n_0_77), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_120 (.ZN (n_0_76), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_119 (.ZN (v[49]), .A1 (n_0_77), .A2 (n_0_76));
NAND2_X1 i_0_118 (.ZN (n_0_75), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_117 (.ZN (n_0_74), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_116 (.ZN (v[48]), .A1 (n_0_75), .A2 (n_0_74));
NAND2_X1 i_0_115 (.ZN (n_0_73), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_114 (.ZN (n_0_72), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_113 (.ZN (v[47]), .A1 (n_0_73), .A2 (n_0_72));
NAND2_X1 i_0_112 (.ZN (n_0_71), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_111 (.ZN (n_0_70), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_110 (.ZN (v[46]), .A1 (n_0_71), .A2 (n_0_70));
NAND2_X1 i_0_109 (.ZN (n_0_69), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_108 (.ZN (n_0_68), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_107 (.ZN (v[45]), .A1 (n_0_69), .A2 (n_0_68));
NAND2_X1 i_0_106 (.ZN (n_0_67), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_105 (.ZN (n_0_66), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_104 (.ZN (v[44]), .A1 (n_0_67), .A2 (n_0_66));
NAND2_X1 i_0_103 (.ZN (n_0_65), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_102 (.ZN (n_0_64), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_101 (.ZN (v[43]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_100 (.ZN (n_0_63), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_99 (.ZN (n_0_62), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_98 (.ZN (v[42]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_97 (.ZN (n_0_61), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_96 (.ZN (n_0_60), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_95 (.ZN (v[41]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_94 (.ZN (n_0_59), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_93 (.ZN (n_0_58), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_92 (.ZN (v[40]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_91 (.ZN (n_0_57), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_90 (.ZN (n_0_56), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_89 (.ZN (v[39]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_88 (.ZN (n_0_55), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_87 (.ZN (n_0_54), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_86 (.ZN (v[38]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_85 (.ZN (n_0_53), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_84 (.ZN (n_0_52), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_83 (.ZN (v[37]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_82 (.ZN (n_0_51), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_81 (.ZN (n_0_50), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_80 (.ZN (v[36]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_79 (.ZN (n_0_49), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_78 (.ZN (n_0_48), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_77 (.ZN (v[35]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_76 (.ZN (n_0_47), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_75 (.ZN (n_0_46), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_74 (.ZN (v[34]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_73 (.ZN (n_0_45), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_72 (.ZN (n_0_44), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_71 (.ZN (v[33]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_70 (.ZN (n_0_43), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_69 (.ZN (n_0_42), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_68 (.ZN (v[32]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_67 (.ZN (n_0_41), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_66 (.ZN (n_0_40), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_65 (.ZN (v[31]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_64 (.ZN (n_0_39), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_63 (.ZN (n_0_38), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_62 (.ZN (v[30]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_61 (.ZN (n_0_37), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_60 (.ZN (n_0_36), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_59 (.ZN (v[29]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_58 (.ZN (n_0_35), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_57 (.ZN (n_0_34), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_56 (.ZN (v[28]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_55 (.ZN (n_0_33), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_54 (.ZN (n_0_32), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_53 (.ZN (v[27]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_52 (.ZN (n_0_31), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_51 (.ZN (n_0_30), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_50 (.ZN (v[26]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_49 (.ZN (n_0_29), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_48 (.ZN (n_0_28), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_47 (.ZN (v[25]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_46 (.ZN (n_0_27), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_45 (.ZN (n_0_26), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_44 (.ZN (v[24]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_43 (.ZN (n_0_25), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_42 (.ZN (n_0_24), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_41 (.ZN (v[23]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_40 (.ZN (n_0_23), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_39 (.ZN (n_0_22), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_38 (.ZN (v[22]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_37 (.ZN (n_0_21), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_36 (.ZN (n_0_20), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_35 (.ZN (v[21]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_34 (.ZN (n_0_19), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_33 (.ZN (n_0_18), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_32 (.ZN (v[20]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_31 (.ZN (n_0_17), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_30 (.ZN (n_0_16), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_29 (.ZN (v[19]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_28 (.ZN (n_0_15), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_27 (.ZN (n_0_14), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_26 (.ZN (v[18]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_25 (.ZN (n_0_13), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_24 (.ZN (n_0_12), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_23 (.ZN (v[17]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_22 (.ZN (n_0_11), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_21 (.ZN (n_0_10), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_20 (.ZN (v[16]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_19 (.ZN (n_0_9), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_18 (.ZN (n_0_8), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_17 (.ZN (v[15]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_16 (.ZN (n_0_7), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_15 (.ZN (n_0_6), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X2 i_0_14 (.ZN (v[14]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_13 (.ZN (n_0_5), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_12 (.ZN (n_0_4), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X2 i_0_11 (.ZN (v[13]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_10 (.ZN (n_0_3), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_9 (.ZN (n_0_2), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X2 i_0_8 (.ZN (v[12]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_7 (.ZN (n_0_1), .A1 (z[10]), .A2 (x[10]));
OAI21_X1 i_0_6 (.ZN (n_0_0), .A (y[10]), .B1 (z[10]), .B2 (x[10]));
NAND2_X1 i_0_5 (.ZN (v[11]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X2 i_0_4 (.ZN (v[10]), .A1 (y[9]), .A2 (x[9]));
AND2_X2 i_0_3 (.ZN (v[9]), .A1 (y[8]), .A2 (x[8]));
AND2_X2 i_0_2 (.ZN (v[8]), .A1 (y[7]), .A2 (x[7]));
AND2_X1 i_0_1 (.ZN (v[7]), .A1 (y[6]), .A2 (x[6]));
AND2_X2 i_0_0 (.ZN (v[6]), .A1 (y[5]), .A2 (x[5]));
XNOR2_X2 slo__mro_c6 (.ZN (slo__mro_n7), .A (y[13]), .B (z[13]));
XNOR2_X2 slo__mro_c7 (.ZN (u[13]), .A (slo__mro_n7), .B (x[13]));

endmodule //CSA__0_75

module CSA__3_14 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_71;
wire n_0_72;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;


INV_X1 i_0_173 (.ZN (n_0_107), .A (y[11]));
INV_X1 i_0_172 (.ZN (n_0_106), .A (x[11]));
NAND2_X1 i_0_171 (.ZN (n_0_105), .A1 (n_0_106), .A2 (z[11]));
INV_X1 i_0_170 (.ZN (n_0_104), .A (z[11]));
NAND2_X1 i_0_169 (.ZN (n_0_103), .A1 (n_0_104), .A2 (x[11]));
NAND2_X1 i_0_168 (.ZN (n_0_102), .A1 (n_0_103), .A2 (n_0_105));
NAND2_X1 i_0_167 (.ZN (n_0_101), .A1 (n_0_102), .A2 (n_0_107));
NAND3_X1 i_0_166 (.ZN (n_0_100), .A1 (n_0_103), .A2 (n_0_105), .A3 (y[11]));
NAND2_X1 i_0_165 (.ZN (u[11]), .A1 (n_0_101), .A2 (n_0_100));
INV_X1 i_0_164 (.ZN (n_0_99), .A (y[10]));
INV_X1 i_0_163 (.ZN (n_0_98), .A (x[10]));
NAND2_X2 i_0_162 (.ZN (n_0_97), .A1 (n_0_98), .A2 (z[10]));
INV_X2 i_0_161 (.ZN (n_0_96), .A (z[10]));
NAND2_X2 i_0_160 (.ZN (n_0_95), .A1 (n_0_96), .A2 (x[10]));
NAND2_X1 i_0_116 (.ZN (n_0_94), .A1 (n_0_95), .A2 (n_0_97));
NAND2_X1 i_0_115 (.ZN (n_0_72), .A1 (n_0_94), .A2 (n_0_99));
NAND3_X1 i_0_114 (.ZN (n_0_71), .A1 (n_0_95), .A2 (n_0_97), .A3 (y[10]));
NAND2_X2 i_0_113 (.ZN (u[10]), .A1 (n_0_71), .A2 (n_0_72));
XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[61]), .B (x[61]));
XOR2_X1 i_0_158 (.Z (u[61]), .A (z[61]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[32]), .A (z[32]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[31]), .B (x[61]));
XNOR2_X1 i_0_155 (.ZN (u[31]), .A (y[31]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_153 (.ZN (u[30]), .A (y[30]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_151 (.ZN (u[29]), .A (y[29]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_149 (.ZN (u[28]), .A (y[28]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_147 (.ZN (u[27]), .A (y[27]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_145 (.ZN (u[26]), .A (y[26]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_143 (.ZN (u[25]), .A (y[25]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_141 (.ZN (u[24]), .A (y[24]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_139 (.ZN (u[23]), .A (y[23]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_137 (.ZN (u[22]), .A (y[22]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_135 (.ZN (u[21]), .A (y[21]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_133 (.ZN (u[20]), .A (y[20]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_131 (.ZN (u[19]), .A (y[19]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_129 (.ZN (u[18]), .A (y[18]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_127 (.ZN (u[17]), .A (y[17]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_125 (.ZN (u[16]), .A (y[16]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[15]), .B (x[15]));
XNOR2_X1 i_0_123 (.ZN (u[15]), .A (y[15]), .B (n_0_76));
XNOR2_X2 i_0_122 (.ZN (n_0_75), .A (z[14]), .B (x[14]));
XNOR2_X1 i_0_121 (.ZN (u[14]), .A (y[14]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[13]), .B (x[13]));
XNOR2_X1 i_0_119 (.ZN (u[13]), .A (y[13]), .B (n_0_74));
XNOR2_X2 i_0_118 (.ZN (n_0_73), .A (z[12]), .B (x[12]));
XNOR2_X2 i_0_117 (.ZN (u[12]), .A (y[12]), .B (n_0_73));
XNOR2_X2 i_0_112 (.ZN (n_0_70), .A (x[9]), .B (z[9]));
XNOR2_X2 i_0_111 (.ZN (u[9]), .A (n_0_70), .B (y[9]));
XNOR2_X2 i_0_110 (.ZN (n_0_69), .A (z[8]), .B (x[8]));
XNOR2_X2 i_0_109 (.ZN (u[8]), .A (y[8]), .B (n_0_69));
XNOR2_X1 i_0_108 (.ZN (n_0_68), .A (z[7]), .B (x[7]));
XNOR2_X1 i_0_107 (.ZN (u[7]), .A (y[7]), .B (n_0_68));
XNOR2_X2 i_0_106 (.ZN (n_0_67), .A (x[6]), .B (z[6]));
XNOR2_X2 i_0_105 (.ZN (u[6]), .A (n_0_67), .B (y[6]));
XNOR2_X1 i_0_104 (.ZN (n_0_66), .A (z[5]), .B (x[5]));
XNOR2_X2 i_0_103 (.ZN (u[5]), .A (y[5]), .B (n_0_66));
XNOR2_X1 i_0_102 (.ZN (n_0_65), .A (z[4]), .B (x[4]));
XNOR2_X1 i_0_101 (.ZN (u[4]), .A (y[4]), .B (n_0_65));
XNOR2_X1 i_0_100 (.ZN (n_0_64), .A (z[3]), .B (x[3]));
XNOR2_X1 i_0_99 (.ZN (u[3]), .A (y[3]), .B (n_0_64));
XNOR2_X1 i_0_98 (.ZN (n_0_63), .A (z[2]), .B (x[2]));
XNOR2_X1 i_0_97 (.ZN (u[2]), .A (y[2]), .B (n_0_63));
XOR2_X1 i_0_96 (.Z (u[1]), .A (y[1]), .B (x[1]));
NAND2_X1 i_0_95 (.ZN (n_0_62), .A1 (y[61]), .A2 (x[61]));
OAI21_X1 i_0_94 (.ZN (n_0_61), .A (z[61]), .B1 (x[61]), .B2 (y[61]));
NAND2_X1 i_0_93 (.ZN (v[61]), .A1 (n_0_62), .A2 (n_0_61));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (z[32]), .B1 (x[61]), .B2 (y[61]));
NAND2_X1 i_0_91 (.ZN (v[33]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[31]), .A2 (x[61]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[31]), .B1 (z[31]), .B2 (x[61]));
NAND2_X1 i_0_88 (.ZN (v[32]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_85 (.ZN (v[31]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_82 (.ZN (v[30]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_79 (.ZN (v[29]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_76 (.ZN (v[28]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_73 (.ZN (v[27]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_70 (.ZN (v[26]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_67 (.ZN (v[25]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_64 (.ZN (v[24]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_61 (.ZN (v[23]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_58 (.ZN (v[22]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_55 (.ZN (v[21]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_52 (.ZN (v[20]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_49 (.ZN (v[19]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_46 (.ZN (v[18]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_43 (.ZN (v[17]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_40 (.ZN (v[16]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_37 (.ZN (v[15]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X1 i_0_34 (.ZN (v[14]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X1 i_0_31 (.ZN (v[13]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X1 i_0_28 (.ZN (v[12]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[10]), .A2 (x[10]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[10]), .B1 (z[10]), .B2 (x[10]));
NAND2_X1 i_0_25 (.ZN (v[11]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[9]), .A2 (x[9]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[9]), .B1 (z[9]), .B2 (x[9]));
NAND2_X2 i_0_22 (.ZN (v[10]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[8]), .A2 (x[8]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[8]), .B1 (z[8]), .B2 (x[8]));
NAND2_X1 i_0_19 (.ZN (v[9]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[7]), .A2 (x[7]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[7]), .B1 (z[7]), .B2 (x[7]));
NAND2_X1 i_0_16 (.ZN (v[8]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[6]), .A2 (x[6]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[6]), .B1 (z[6]), .B2 (x[6]));
NAND2_X1 i_0_13 (.ZN (v[7]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[5]), .A2 (x[5]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[5]), .B1 (z[5]), .B2 (x[5]));
NAND2_X1 i_0_10 (.ZN (v[6]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[4]), .A2 (x[4]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[4]), .B1 (z[4]), .B2 (x[4]));
NAND2_X1 i_0_7 (.ZN (v[5]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[3]), .A2 (x[3]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[3]), .B1 (z[3]), .B2 (x[3]));
NAND2_X1 i_0_4 (.ZN (v[4]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[2]), .A2 (x[2]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[2]), .B1 (z[2]), .B2 (x[2]));
NAND2_X1 i_0_1 (.ZN (v[3]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[2]), .A1 (y[1]), .A2 (x[1]));

endmodule //CSA__3_14

module CSA__3_11 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire slo__sro_n39;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire slo__sro_n30;
wire n_0_66;
wire n_0_67;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_69;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_8;
wire n_0_68;
wire slo__mro_n15;


NAND2_X1 i_0_172 (.ZN (n_0_68), .A1 (y[9]), .A2 (x[9]));
NAND2_X2 i_0_170 (.ZN (v[10]), .A1 (slo__sro_n39), .A2 (n_0_68));
INV_X1 i_0_174 (.ZN (n_0_8), .A (y[11]));
INV_X1 i_0_169 (.ZN (n_0_107), .A (x[11]));
NAND2_X1 i_0_167 (.ZN (n_0_106), .A1 (n_0_107), .A2 (z[11]));
INV_X1 i_0_107 (.ZN (n_0_105), .A (z[11]));
NAND2_X2 i_0_15 (.ZN (n_0_104), .A1 (n_0_105), .A2 (x[11]));
NAND2_X1 i_0_14 (.ZN (n_0_103), .A1 (n_0_106), .A2 (n_0_104));
NAND2_X1 i_0_168 (.ZN (n_0_102), .A1 (n_0_103), .A2 (n_0_8));
NAND3_X2 i_0_13 (.ZN (n_0_101), .A1 (n_0_106), .A2 (n_0_104), .A3 (y[11]));
NAND2_X2 i_0_166 (.ZN (u[11]), .A1 (n_0_102), .A2 (n_0_101));
INV_X1 i_0_165 (.ZN (n_0_100), .A (y[10]));
INV_X2 i_0_164 (.ZN (n_0_99), .A (x[10]));
NAND2_X2 i_0_163 (.ZN (n_0_98), .A1 (n_0_99), .A2 (z[10]));
INV_X2 i_0_162 (.ZN (n_0_97), .A (z[10]));
NAND2_X2 i_0_161 (.ZN (n_0_96), .A1 (n_0_97), .A2 (x[10]));
NAND2_X1 i_0_160 (.ZN (n_0_95), .A1 (n_0_98), .A2 (n_0_96));
NAND3_X1 i_0_109 (.ZN (n_0_69), .A1 (n_0_96), .A2 (n_0_98), .A3 (y[10]));
NAND2_X2 i_0_108 (.ZN (u[10]), .A1 (n_0_69), .A2 (slo__sro_n30));
XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[62]), .B (x[62]));
XOR2_X1 i_0_158 (.Z (u[61]), .A (z[62]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[35]), .A (z[35]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[34]), .B (x[62]));
XNOR2_X1 i_0_155 (.ZN (u[34]), .A (y[34]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_153 (.ZN (u[33]), .A (y[33]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_151 (.ZN (u[32]), .A (y[32]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_149 (.ZN (u[31]), .A (y[31]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_147 (.ZN (u[30]), .A (y[30]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_145 (.ZN (u[29]), .A (y[29]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_143 (.ZN (u[28]), .A (y[28]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_141 (.ZN (u[27]), .A (y[27]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_139 (.ZN (u[26]), .A (y[26]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_137 (.ZN (u[25]), .A (y[25]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_135 (.ZN (u[24]), .A (y[24]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_133 (.ZN (u[23]), .A (y[23]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_131 (.ZN (u[22]), .A (y[22]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_129 (.ZN (u[21]), .A (y[21]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_127 (.ZN (u[20]), .A (y[20]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_125 (.ZN (u[19]), .A (y[19]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_123 (.ZN (u[18]), .A (y[18]), .B (n_0_76));
XNOR2_X1 i_0_122 (.ZN (n_0_75), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_121 (.ZN (u[17]), .A (y[17]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_119 (.ZN (u[16]), .A (y[16]), .B (n_0_74));
XNOR2_X1 i_0_118 (.ZN (n_0_73), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_117 (.ZN (u[15]), .A (y[15]), .B (n_0_73));
XNOR2_X1 i_0_116 (.ZN (n_0_72), .A (z[14]), .B (x[14]));
XNOR2_X1 i_0_115 (.ZN (u[14]), .A (y[14]), .B (n_0_72));
XNOR2_X2 i_0_114 (.ZN (n_0_71), .A (z[13]), .B (x[13]));
XNOR2_X2 i_0_113 (.ZN (u[13]), .A (y[13]), .B (n_0_71));
XNOR2_X2 i_0_112 (.ZN (n_0_70), .A (z[12]), .B (x[12]));
XNOR2_X2 i_0_111 (.ZN (u[12]), .A (n_0_70), .B (y[12]));
XNOR2_X1 i_0_106 (.ZN (n_0_67), .A (x[9]), .B (z[9]));
XNOR2_X2 i_0_105 (.ZN (u[9]), .A (n_0_67), .B (y[9]));
XNOR2_X2 i_0_104 (.ZN (n_0_66), .A (z[8]), .B (x[8]));
XNOR2_X2 i_0_103 (.ZN (u[8]), .A (n_0_66), .B (y[8]));
NAND2_X2 slo__sro_c42 (.ZN (slo__sro_n30), .A1 (n_0_95), .A2 (n_0_100));
OAI21_X1 slo__sro_c51 (.ZN (slo__sro_n39), .A (z[9]), .B1 (x[9]), .B2 (y[9]));
XNOR2_X1 i_0_100 (.ZN (n_0_64), .A (z[6]), .B (x[6]));
XNOR2_X2 i_0_99 (.ZN (u[6]), .A (y[6]), .B (n_0_64));
XNOR2_X2 i_0_98 (.ZN (n_0_63), .A (z[5]), .B (x[5]));
XNOR2_X2 i_0_97 (.ZN (u[5]), .A (y[5]), .B (n_0_63));
XOR2_X1 i_0_96 (.Z (u[4]), .A (y[4]), .B (x[4]));
NAND2_X2 i_0_95 (.ZN (n_0_62), .A1 (y[62]), .A2 (x[62]));
OAI21_X1 i_0_94 (.ZN (n_0_61), .A (z[62]), .B1 (x[62]), .B2 (y[62]));
NAND2_X4 i_0_93 (.ZN (v[63]), .A1 (n_0_62), .A2 (n_0_61));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (z[35]), .B1 (x[62]), .B2 (y[62]));
NAND2_X1 i_0_91 (.ZN (v[36]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[34]), .A2 (x[62]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[34]), .B1 (z[34]), .B2 (x[62]));
NAND2_X1 i_0_88 (.ZN (v[35]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_85 (.ZN (v[34]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_82 (.ZN (v[33]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_79 (.ZN (v[32]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_76 (.ZN (v[31]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_73 (.ZN (v[30]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_70 (.ZN (v[29]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_67 (.ZN (v[28]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_64 (.ZN (v[27]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_61 (.ZN (v[26]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_58 (.ZN (v[25]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_55 (.ZN (v[24]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_52 (.ZN (v[23]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_49 (.ZN (v[22]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_46 (.ZN (v[21]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_43 (.ZN (v[20]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_40 (.ZN (v[19]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_37 (.ZN (v[18]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_34 (.ZN (v[17]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_31 (.ZN (v[16]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_28 (.ZN (v[15]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X1 i_0_25 (.ZN (v[14]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X2 i_0_22 (.ZN (v[13]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X1 i_0_19 (.ZN (v[12]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[10]), .A2 (x[10]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[10]), .B1 (z[10]), .B2 (x[10]));
NAND2_X1 i_0_16 (.ZN (v[11]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[8]), .A2 (x[8]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[8]), .B1 (z[8]), .B2 (x[8]));
NAND2_X2 i_0_10 (.ZN (v[9]), .A1 (n_0_6), .A2 (n_0_7));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[7]), .A2 (x[7]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[7]), .B1 (z[7]), .B2 (x[7]));
NAND2_X2 i_0_7 (.ZN (v[8]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[6]), .A2 (x[6]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[6]), .B1 (z[6]), .B2 (x[6]));
NAND2_X1 i_0_4 (.ZN (v[7]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[5]), .A2 (x[5]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[5]), .B1 (z[5]), .B2 (x[5]));
NAND2_X1 i_0_1 (.ZN (v[6]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[5]), .A1 (y[4]), .A2 (x[4]));
XNOR2_X2 slo__mro_c28 (.ZN (slo__mro_n15), .A (x[7]), .B (z[7]));
XNOR2_X2 slo__mro_c29 (.ZN (u[7]), .A (slo__mro_n15), .B (y[7]));

endmodule //CSA__3_11

module CSA__3_8 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire slo__mro_n51;
wire slo__mro_n16;
wire n_0_0;
wire n_0_1;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire slo__mro_n3;


XNOR2_X1 i_0_287 (.ZN (n_0_168), .A (z[63]), .B (x[63]));
XNOR2_X1 i_0_286 (.ZN (u[63]), .A (y[63]), .B (n_0_168));
XNOR2_X1 i_0_285 (.ZN (n_0_167), .A (z[62]), .B (x[62]));
XNOR2_X1 i_0_284 (.ZN (u[62]), .A (y[62]), .B (n_0_167));
XNOR2_X1 i_0_283 (.ZN (n_0_166), .A (z[61]), .B (x[61]));
XNOR2_X1 i_0_282 (.ZN (u[61]), .A (y[61]), .B (n_0_166));
XNOR2_X1 i_0_281 (.ZN (n_0_165), .A (z[60]), .B (x[60]));
XNOR2_X1 i_0_280 (.ZN (u[60]), .A (y[60]), .B (n_0_165));
XNOR2_X1 i_0_279 (.ZN (n_0_164), .A (z[59]), .B (x[59]));
XNOR2_X1 i_0_278 (.ZN (u[59]), .A (y[59]), .B (n_0_164));
XNOR2_X1 i_0_277 (.ZN (n_0_163), .A (z[58]), .B (x[58]));
XNOR2_X1 i_0_276 (.ZN (u[58]), .A (y[58]), .B (n_0_163));
XNOR2_X1 i_0_275 (.ZN (n_0_162), .A (z[57]), .B (x[57]));
XNOR2_X1 i_0_274 (.ZN (u[57]), .A (y[57]), .B (n_0_162));
XNOR2_X1 i_0_273 (.ZN (n_0_161), .A (z[56]), .B (x[56]));
XNOR2_X1 i_0_272 (.ZN (u[56]), .A (y[56]), .B (n_0_161));
XNOR2_X1 i_0_271 (.ZN (n_0_160), .A (z[55]), .B (x[55]));
XNOR2_X1 i_0_270 (.ZN (u[55]), .A (y[55]), .B (n_0_160));
XNOR2_X1 i_0_269 (.ZN (n_0_159), .A (z[54]), .B (x[54]));
XNOR2_X1 i_0_268 (.ZN (u[54]), .A (y[54]), .B (n_0_159));
XNOR2_X1 i_0_267 (.ZN (n_0_158), .A (z[53]), .B (x[53]));
XNOR2_X1 i_0_266 (.ZN (u[53]), .A (y[53]), .B (n_0_158));
XNOR2_X1 i_0_265 (.ZN (n_0_157), .A (z[52]), .B (x[52]));
XNOR2_X1 i_0_264 (.ZN (u[52]), .A (y[52]), .B (n_0_157));
XNOR2_X1 i_0_263 (.ZN (n_0_156), .A (z[51]), .B (x[51]));
XNOR2_X1 i_0_262 (.ZN (u[51]), .A (y[51]), .B (n_0_156));
XNOR2_X1 i_0_261 (.ZN (n_0_155), .A (z[50]), .B (x[50]));
XNOR2_X1 i_0_260 (.ZN (u[50]), .A (y[50]), .B (n_0_155));
XNOR2_X1 i_0_259 (.ZN (n_0_154), .A (z[49]), .B (x[49]));
XNOR2_X1 i_0_258 (.ZN (u[49]), .A (y[49]), .B (n_0_154));
XNOR2_X1 i_0_257 (.ZN (n_0_153), .A (z[48]), .B (x[48]));
XNOR2_X1 i_0_256 (.ZN (u[48]), .A (y[48]), .B (n_0_153));
XNOR2_X1 i_0_255 (.ZN (n_0_152), .A (z[47]), .B (x[47]));
XNOR2_X1 i_0_254 (.ZN (u[47]), .A (y[47]), .B (n_0_152));
XNOR2_X1 i_0_253 (.ZN (n_0_151), .A (z[46]), .B (x[46]));
XNOR2_X1 i_0_252 (.ZN (u[46]), .A (y[46]), .B (n_0_151));
XNOR2_X1 i_0_251 (.ZN (n_0_150), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_250 (.ZN (u[45]), .A (y[45]), .B (n_0_150));
XNOR2_X1 i_0_249 (.ZN (n_0_149), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_248 (.ZN (u[44]), .A (y[44]), .B (n_0_149));
XNOR2_X1 i_0_247 (.ZN (n_0_148), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_246 (.ZN (u[43]), .A (y[43]), .B (n_0_148));
XNOR2_X1 i_0_245 (.ZN (n_0_147), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_244 (.ZN (u[42]), .A (y[42]), .B (n_0_147));
XNOR2_X1 i_0_243 (.ZN (n_0_146), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_242 (.ZN (u[41]), .A (y[41]), .B (n_0_146));
XNOR2_X1 i_0_241 (.ZN (n_0_145), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_240 (.ZN (u[40]), .A (y[40]), .B (n_0_145));
XNOR2_X1 i_0_239 (.ZN (n_0_144), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_238 (.ZN (u[39]), .A (y[39]), .B (n_0_144));
XNOR2_X1 i_0_237 (.ZN (n_0_143), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_236 (.ZN (u[38]), .A (y[38]), .B (n_0_143));
XNOR2_X1 i_0_235 (.ZN (n_0_142), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_234 (.ZN (u[37]), .A (y[37]), .B (n_0_142));
XNOR2_X1 i_0_233 (.ZN (n_0_141), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_232 (.ZN (u[36]), .A (y[36]), .B (n_0_141));
XNOR2_X1 i_0_231 (.ZN (n_0_140), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_230 (.ZN (u[35]), .A (y[35]), .B (n_0_140));
XNOR2_X1 i_0_229 (.ZN (n_0_139), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_228 (.ZN (u[34]), .A (y[34]), .B (n_0_139));
XNOR2_X1 i_0_227 (.ZN (n_0_138), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_226 (.ZN (u[33]), .A (y[33]), .B (n_0_138));
XNOR2_X1 i_0_225 (.ZN (n_0_137), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_224 (.ZN (u[32]), .A (y[32]), .B (n_0_137));
XNOR2_X1 i_0_223 (.ZN (n_0_136), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_222 (.ZN (u[31]), .A (y[31]), .B (n_0_136));
XNOR2_X1 i_0_221 (.ZN (n_0_135), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_220 (.ZN (u[30]), .A (y[30]), .B (n_0_135));
XNOR2_X1 i_0_219 (.ZN (n_0_134), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_218 (.ZN (u[29]), .A (y[29]), .B (n_0_134));
XNOR2_X1 i_0_217 (.ZN (n_0_133), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_216 (.ZN (u[28]), .A (y[28]), .B (n_0_133));
XNOR2_X1 i_0_215 (.ZN (n_0_132), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_214 (.ZN (u[27]), .A (y[27]), .B (n_0_132));
XNOR2_X1 i_0_213 (.ZN (n_0_131), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_212 (.ZN (u[26]), .A (y[26]), .B (n_0_131));
XNOR2_X1 i_0_211 (.ZN (n_0_130), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_210 (.ZN (u[25]), .A (y[25]), .B (n_0_130));
XNOR2_X1 i_0_209 (.ZN (n_0_129), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_208 (.ZN (u[24]), .A (y[24]), .B (n_0_129));
XNOR2_X1 i_0_207 (.ZN (n_0_128), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_206 (.ZN (u[23]), .A (y[23]), .B (n_0_128));
XNOR2_X1 i_0_205 (.ZN (n_0_127), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_204 (.ZN (u[22]), .A (y[22]), .B (n_0_127));
XNOR2_X1 i_0_203 (.ZN (n_0_126), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_202 (.ZN (u[21]), .A (y[21]), .B (n_0_126));
XNOR2_X1 i_0_201 (.ZN (n_0_125), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_200 (.ZN (u[20]), .A (y[20]), .B (n_0_125));
XNOR2_X1 i_0_199 (.ZN (n_0_124), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_198 (.ZN (u[19]), .A (y[19]), .B (n_0_124));
XNOR2_X1 i_0_197 (.ZN (n_0_123), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_196 (.ZN (u[18]), .A (y[18]), .B (n_0_123));
XNOR2_X1 i_0_195 (.ZN (n_0_122), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_194 (.ZN (u[17]), .A (y[17]), .B (n_0_122));
XNOR2_X2 i_0_193 (.ZN (n_0_121), .A (z[16]), .B (x[16]));
XNOR2_X2 i_0_192 (.ZN (u[16]), .A (y[16]), .B (n_0_121));
XNOR2_X2 i_0_191 (.ZN (n_0_120), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_190 (.ZN (u[15]), .A (n_0_120), .B (y[15]));
XNOR2_X2 i_0_189 (.ZN (n_0_119), .A (z[14]), .B (x[14]));
XNOR2_X2 i_0_188 (.ZN (u[14]), .A (y[14]), .B (n_0_119));
XNOR2_X2 i_0_187 (.ZN (n_0_118), .A (z[13]), .B (x[13]));
XNOR2_X2 i_0_186 (.ZN (u[13]), .A (y[13]), .B (n_0_118));
XNOR2_X2 i_0_185 (.ZN (n_0_117), .A (z[12]), .B (x[12]));
XNOR2_X2 i_0_184 (.ZN (u[12]), .A (n_0_117), .B (y[12]));
XNOR2_X2 i_0_183 (.ZN (n_0_116), .A (x[11]), .B (z[11]));
XNOR2_X2 i_0_182 (.ZN (u[11]), .A (n_0_116), .B (y[11]));
XNOR2_X2 i_0_181 (.ZN (n_0_115), .A (x[10]), .B (z[10]));
XNOR2_X2 i_0_180 (.ZN (u[10]), .A (n_0_115), .B (y[10]));
XNOR2_X2 i_0_179 (.ZN (n_0_114), .A (x[9]), .B (z[9]));
XNOR2_X2 i_0_178 (.ZN (u[9]), .A (n_0_114), .B (y[9]));
OAI21_X1 slo__mro_c38 (.ZN (slo__mro_n51), .A (y[8]), .B1 (x[8]), .B2 (z[8]));
NAND2_X1 slo__mro_c39 (.ZN (v[9]), .A1 (slo__mro_n51), .A2 (n_0_3));
XNOR2_X2 slo__mro_c12 (.ZN (slo__mro_n16), .A (y[8]), .B (z[8]));
XNOR2_X2 slo__mro_c13 (.ZN (u[8]), .A (slo__mro_n16), .B (x[8]));
XOR2_X2 i_0_173 (.Z (u[6]), .A (y[6]), .B (x[6]));
XOR2_X1 i_0_172 (.Z (u[5]), .A (y[5]), .B (x[5]));
XOR2_X1 i_0_171 (.Z (u[4]), .A (y[4]), .B (x[4]));
NAND2_X1 i_0_170 (.ZN (n_0_111), .A1 (z[62]), .A2 (x[62]));
OAI21_X1 i_0_169 (.ZN (n_0_110), .A (y[62]), .B1 (z[62]), .B2 (x[62]));
NAND2_X1 i_0_168 (.ZN (v[63]), .A1 (n_0_111), .A2 (n_0_110));
NAND2_X1 i_0_167 (.ZN (n_0_109), .A1 (z[61]), .A2 (x[61]));
OAI21_X1 i_0_166 (.ZN (n_0_108), .A (y[61]), .B1 (z[61]), .B2 (x[61]));
NAND2_X1 i_0_165 (.ZN (v[62]), .A1 (n_0_109), .A2 (n_0_108));
NAND2_X1 i_0_164 (.ZN (n_0_107), .A1 (z[60]), .A2 (x[60]));
OAI21_X1 i_0_163 (.ZN (n_0_106), .A (y[60]), .B1 (z[60]), .B2 (x[60]));
NAND2_X1 i_0_162 (.ZN (v[61]), .A1 (n_0_107), .A2 (n_0_106));
NAND2_X1 i_0_161 (.ZN (n_0_105), .A1 (z[59]), .A2 (x[59]));
OAI21_X1 i_0_160 (.ZN (n_0_104), .A (y[59]), .B1 (z[59]), .B2 (x[59]));
NAND2_X1 i_0_159 (.ZN (v[60]), .A1 (n_0_105), .A2 (n_0_104));
NAND2_X1 i_0_158 (.ZN (n_0_103), .A1 (z[58]), .A2 (x[58]));
OAI21_X1 i_0_157 (.ZN (n_0_102), .A (y[58]), .B1 (z[58]), .B2 (x[58]));
NAND2_X1 i_0_156 (.ZN (v[59]), .A1 (n_0_103), .A2 (n_0_102));
NAND2_X1 i_0_155 (.ZN (n_0_101), .A1 (z[57]), .A2 (x[57]));
OAI21_X1 i_0_154 (.ZN (n_0_100), .A (y[57]), .B1 (z[57]), .B2 (x[57]));
NAND2_X1 i_0_153 (.ZN (v[58]), .A1 (n_0_101), .A2 (n_0_100));
NAND2_X1 i_0_152 (.ZN (n_0_99), .A1 (z[56]), .A2 (x[56]));
OAI21_X1 i_0_151 (.ZN (n_0_98), .A (y[56]), .B1 (z[56]), .B2 (x[56]));
NAND2_X1 i_0_150 (.ZN (v[57]), .A1 (n_0_99), .A2 (n_0_98));
NAND2_X1 i_0_149 (.ZN (n_0_97), .A1 (z[55]), .A2 (x[55]));
OAI21_X1 i_0_148 (.ZN (n_0_96), .A (y[55]), .B1 (z[55]), .B2 (x[55]));
NAND2_X1 i_0_147 (.ZN (v[56]), .A1 (n_0_97), .A2 (n_0_96));
NAND2_X1 i_0_146 (.ZN (n_0_95), .A1 (z[54]), .A2 (x[54]));
OAI21_X1 i_0_145 (.ZN (n_0_94), .A (y[54]), .B1 (z[54]), .B2 (x[54]));
NAND2_X1 i_0_144 (.ZN (v[55]), .A1 (n_0_95), .A2 (n_0_94));
NAND2_X1 i_0_143 (.ZN (n_0_93), .A1 (z[53]), .A2 (x[53]));
OAI21_X1 i_0_142 (.ZN (n_0_92), .A (y[53]), .B1 (z[53]), .B2 (x[53]));
NAND2_X1 i_0_141 (.ZN (v[54]), .A1 (n_0_93), .A2 (n_0_92));
NAND2_X1 i_0_140 (.ZN (n_0_91), .A1 (z[52]), .A2 (x[52]));
OAI21_X1 i_0_139 (.ZN (n_0_90), .A (y[52]), .B1 (z[52]), .B2 (x[52]));
NAND2_X1 i_0_138 (.ZN (v[53]), .A1 (n_0_91), .A2 (n_0_90));
NAND2_X1 i_0_137 (.ZN (n_0_89), .A1 (z[51]), .A2 (x[51]));
OAI21_X1 i_0_136 (.ZN (n_0_88), .A (y[51]), .B1 (z[51]), .B2 (x[51]));
NAND2_X1 i_0_135 (.ZN (v[52]), .A1 (n_0_89), .A2 (n_0_88));
NAND2_X1 i_0_134 (.ZN (n_0_87), .A1 (z[50]), .A2 (x[50]));
OAI21_X1 i_0_133 (.ZN (n_0_86), .A (y[50]), .B1 (z[50]), .B2 (x[50]));
NAND2_X1 i_0_132 (.ZN (v[51]), .A1 (n_0_87), .A2 (n_0_86));
NAND2_X1 i_0_131 (.ZN (n_0_85), .A1 (z[49]), .A2 (x[49]));
OAI21_X1 i_0_130 (.ZN (n_0_84), .A (y[49]), .B1 (z[49]), .B2 (x[49]));
NAND2_X1 i_0_129 (.ZN (v[50]), .A1 (n_0_85), .A2 (n_0_84));
NAND2_X1 i_0_128 (.ZN (n_0_83), .A1 (z[48]), .A2 (x[48]));
OAI21_X1 i_0_127 (.ZN (n_0_82), .A (y[48]), .B1 (z[48]), .B2 (x[48]));
NAND2_X1 i_0_126 (.ZN (v[49]), .A1 (n_0_83), .A2 (n_0_82));
NAND2_X1 i_0_125 (.ZN (n_0_81), .A1 (z[47]), .A2 (x[47]));
OAI21_X1 i_0_124 (.ZN (n_0_80), .A (y[47]), .B1 (z[47]), .B2 (x[47]));
NAND2_X1 i_0_123 (.ZN (v[48]), .A1 (n_0_81), .A2 (n_0_80));
NAND2_X1 i_0_122 (.ZN (n_0_79), .A1 (z[46]), .A2 (x[46]));
OAI21_X1 i_0_121 (.ZN (n_0_78), .A (y[46]), .B1 (z[46]), .B2 (x[46]));
NAND2_X1 i_0_120 (.ZN (v[47]), .A1 (n_0_79), .A2 (n_0_78));
NAND2_X1 i_0_119 (.ZN (n_0_77), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_118 (.ZN (n_0_76), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_117 (.ZN (v[46]), .A1 (n_0_77), .A2 (n_0_76));
NAND2_X1 i_0_116 (.ZN (n_0_75), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_115 (.ZN (n_0_74), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_114 (.ZN (v[45]), .A1 (n_0_75), .A2 (n_0_74));
NAND2_X1 i_0_113 (.ZN (n_0_73), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_112 (.ZN (n_0_72), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_111 (.ZN (v[44]), .A1 (n_0_73), .A2 (n_0_72));
NAND2_X1 i_0_110 (.ZN (n_0_71), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_109 (.ZN (n_0_70), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_108 (.ZN (v[43]), .A1 (n_0_71), .A2 (n_0_70));
NAND2_X1 i_0_107 (.ZN (n_0_69), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_106 (.ZN (n_0_68), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_105 (.ZN (v[42]), .A1 (n_0_69), .A2 (n_0_68));
NAND2_X1 i_0_104 (.ZN (n_0_67), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_103 (.ZN (n_0_66), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_102 (.ZN (v[41]), .A1 (n_0_67), .A2 (n_0_66));
NAND2_X1 i_0_101 (.ZN (n_0_65), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_100 (.ZN (n_0_64), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_99 (.ZN (v[40]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_98 (.ZN (n_0_63), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_97 (.ZN (n_0_62), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_96 (.ZN (v[39]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_95 (.ZN (n_0_61), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_94 (.ZN (n_0_60), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_93 (.ZN (v[38]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_92 (.ZN (n_0_59), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_91 (.ZN (n_0_58), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_90 (.ZN (v[37]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_89 (.ZN (n_0_57), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_88 (.ZN (n_0_56), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_87 (.ZN (v[36]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_86 (.ZN (n_0_55), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_85 (.ZN (n_0_54), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_84 (.ZN (v[35]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_83 (.ZN (n_0_53), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_82 (.ZN (n_0_52), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_81 (.ZN (v[34]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_80 (.ZN (n_0_51), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_79 (.ZN (n_0_50), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_78 (.ZN (v[33]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_77 (.ZN (n_0_49), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_76 (.ZN (n_0_48), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_75 (.ZN (v[32]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_74 (.ZN (n_0_47), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_73 (.ZN (n_0_46), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_72 (.ZN (v[31]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_71 (.ZN (n_0_45), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_70 (.ZN (n_0_44), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_69 (.ZN (v[30]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_68 (.ZN (n_0_43), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_67 (.ZN (n_0_42), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_66 (.ZN (v[29]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_65 (.ZN (n_0_41), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_64 (.ZN (n_0_40), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_63 (.ZN (v[28]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_62 (.ZN (n_0_39), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_61 (.ZN (n_0_38), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_60 (.ZN (v[27]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_59 (.ZN (n_0_37), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_58 (.ZN (n_0_36), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_57 (.ZN (v[26]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_56 (.ZN (n_0_35), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_55 (.ZN (n_0_34), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_54 (.ZN (v[25]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_53 (.ZN (n_0_33), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_52 (.ZN (n_0_32), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_51 (.ZN (v[24]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_50 (.ZN (n_0_31), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_49 (.ZN (n_0_30), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_48 (.ZN (v[23]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_47 (.ZN (n_0_29), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_46 (.ZN (n_0_28), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_45 (.ZN (v[22]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_44 (.ZN (n_0_27), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_43 (.ZN (n_0_26), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_42 (.ZN (v[21]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_41 (.ZN (n_0_25), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_40 (.ZN (n_0_24), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_39 (.ZN (v[20]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_38 (.ZN (n_0_23), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_37 (.ZN (n_0_22), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_36 (.ZN (v[19]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_35 (.ZN (n_0_21), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_34 (.ZN (n_0_20), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_33 (.ZN (v[18]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_32 (.ZN (n_0_19), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_31 (.ZN (n_0_18), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_30 (.ZN (v[17]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_29 (.ZN (n_0_17), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_28 (.ZN (n_0_16), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_27 (.ZN (v[16]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_26 (.ZN (n_0_15), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_25 (.ZN (n_0_14), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X2 i_0_24 (.ZN (v[15]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_23 (.ZN (n_0_13), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_22 (.ZN (n_0_12), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X2 i_0_21 (.ZN (v[14]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_20 (.ZN (n_0_11), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_19 (.ZN (n_0_10), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X2 i_0_18 (.ZN (v[13]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_17 (.ZN (n_0_9), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_16 (.ZN (n_0_8), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X2 i_0_15 (.ZN (v[12]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_14 (.ZN (n_0_7), .A1 (z[10]), .A2 (x[10]));
OAI21_X1 i_0_13 (.ZN (n_0_6), .A (y[10]), .B1 (z[10]), .B2 (x[10]));
NAND2_X1 i_0_12 (.ZN (v[11]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_11 (.ZN (n_0_5), .A1 (z[9]), .A2 (x[9]));
OAI21_X1 i_0_10 (.ZN (n_0_4), .A (y[9]), .B1 (z[9]), .B2 (x[9]));
NAND2_X1 i_0_9 (.ZN (v[10]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_8 (.ZN (n_0_3), .A1 (z[8]), .A2 (x[8]));
NAND2_X1 i_0_5 (.ZN (n_0_1), .A1 (z[7]), .A2 (x[7]));
OAI21_X1 i_0_4 (.ZN (n_0_0), .A (y[7]), .B1 (z[7]), .B2 (x[7]));
NAND2_X2 i_0_3 (.ZN (v[8]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X2 i_0_2 (.ZN (v[7]), .A1 (y[6]), .A2 (x[6]));
AND2_X2 i_0_1 (.ZN (v[6]), .A1 (y[5]), .A2 (x[5]));
AND2_X2 i_0_0 (.ZN (v[5]), .A1 (y[4]), .A2 (x[4]));
XNOR2_X2 slo__mro_c1 (.ZN (slo__mro_n3), .A (x[7]), .B (z[7]));
XNOR2_X2 slo__mro_c2 (.ZN (u[7]), .A (slo__mro_n3), .B (y[7]));

endmodule //CSA__3_8

module CSA__3_5 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire slo__mro_n3;


INV_X1 i_0_168 (.ZN (n_0_98), .A (z[61]));
INV_X1 i_0_167 (.ZN (n_0_97), .A (z[35]));
INV_X1 i_0_166 (.ZN (n_0_96), .A (z[34]));
XOR2_X1 i_0_165 (.Z (n_0_95), .A (y[61]), .B (x[61]));
XNOR2_X1 i_0_164 (.ZN (u[62]), .A (n_0_98), .B (n_0_95));
XNOR2_X1 i_0_163 (.ZN (u[35]), .A (n_0_97), .B (n_0_95));
XNOR2_X1 i_0_162 (.ZN (u[34]), .A (n_0_96), .B (n_0_95));
XNOR2_X1 i_0_161 (.ZN (n_0_94), .A (z[33]), .B (x[61]));
XNOR2_X1 i_0_160 (.ZN (u[33]), .A (y[33]), .B (n_0_94));
XNOR2_X1 i_0_159 (.ZN (n_0_93), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_158 (.ZN (u[32]), .A (y[32]), .B (n_0_93));
XNOR2_X1 i_0_157 (.ZN (n_0_92), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_156 (.ZN (u[31]), .A (y[31]), .B (n_0_92));
XNOR2_X1 i_0_155 (.ZN (n_0_91), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_154 (.ZN (u[30]), .A (y[30]), .B (n_0_91));
XNOR2_X1 i_0_153 (.ZN (n_0_90), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_152 (.ZN (u[29]), .A (y[29]), .B (n_0_90));
XNOR2_X1 i_0_151 (.ZN (n_0_89), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_150 (.ZN (u[28]), .A (y[28]), .B (n_0_89));
XNOR2_X1 i_0_149 (.ZN (n_0_88), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_148 (.ZN (u[27]), .A (y[27]), .B (n_0_88));
XNOR2_X1 i_0_147 (.ZN (n_0_87), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_146 (.ZN (u[26]), .A (y[26]), .B (n_0_87));
XNOR2_X1 i_0_145 (.ZN (n_0_86), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_144 (.ZN (u[25]), .A (y[25]), .B (n_0_86));
XNOR2_X1 i_0_143 (.ZN (n_0_85), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_142 (.ZN (u[24]), .A (y[24]), .B (n_0_85));
XNOR2_X1 i_0_141 (.ZN (n_0_84), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_140 (.ZN (u[23]), .A (y[23]), .B (n_0_84));
XNOR2_X1 i_0_139 (.ZN (n_0_83), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_138 (.ZN (u[22]), .A (y[22]), .B (n_0_83));
XNOR2_X1 i_0_137 (.ZN (n_0_82), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_136 (.ZN (u[21]), .A (y[21]), .B (n_0_82));
XNOR2_X1 i_0_135 (.ZN (n_0_81), .A (z[20]), .B (x[20]));
XNOR2_X2 i_0_134 (.ZN (u[20]), .A (y[20]), .B (n_0_81));
XNOR2_X1 i_0_133 (.ZN (n_0_80), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_132 (.ZN (u[19]), .A (y[19]), .B (n_0_80));
XNOR2_X1 i_0_131 (.ZN (n_0_79), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_130 (.ZN (u[18]), .A (y[18]), .B (n_0_79));
XNOR2_X1 i_0_129 (.ZN (n_0_78), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_128 (.ZN (u[17]), .A (y[17]), .B (n_0_78));
XNOR2_X1 i_0_127 (.ZN (n_0_77), .A (z[16]), .B (x[16]));
XNOR2_X2 i_0_126 (.ZN (u[16]), .A (y[16]), .B (n_0_77));
XNOR2_X2 i_0_125 (.ZN (n_0_76), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_124 (.ZN (u[15]), .A (y[15]), .B (n_0_76));
XNOR2_X2 i_0_123 (.ZN (n_0_75), .A (z[14]), .B (x[14]));
XNOR2_X2 i_0_122 (.ZN (u[14]), .A (y[14]), .B (n_0_75));
XNOR2_X2 i_0_121 (.ZN (n_0_74), .A (z[13]), .B (x[13]));
XNOR2_X2 i_0_120 (.ZN (u[13]), .A (y[13]), .B (n_0_74));
XNOR2_X2 i_0_119 (.ZN (n_0_73), .A (z[12]), .B (x[12]));
XNOR2_X2 i_0_118 (.ZN (u[12]), .A (n_0_73), .B (y[12]));
XNOR2_X2 i_0_117 (.ZN (n_0_72), .A (z[11]), .B (x[11]));
XNOR2_X2 i_0_116 (.ZN (u[11]), .A (n_0_72), .B (y[11]));
XNOR2_X2 i_0_115 (.ZN (n_0_71), .A (z[10]), .B (x[10]));
XNOR2_X2 i_0_114 (.ZN (u[10]), .A (n_0_71), .B (y[10]));
XNOR2_X2 i_0_113 (.ZN (n_0_70), .A (x[9]), .B (z[9]));
XNOR2_X2 i_0_112 (.ZN (u[9]), .A (n_0_70), .B (y[9]));
XNOR2_X2 i_0_111 (.ZN (n_0_69), .A (z[8]), .B (x[8]));
XNOR2_X2 i_0_110 (.ZN (u[8]), .A (n_0_69), .B (y[8]));
XNOR2_X2 i_0_109 (.ZN (n_0_68), .A (z[7]), .B (x[7]));
XNOR2_X2 i_0_108 (.ZN (u[7]), .A (n_0_68), .B (y[7]));
XNOR2_X2 i_0_107 (.ZN (n_0_67), .A (z[6]), .B (x[6]));
XNOR2_X2 i_0_106 (.ZN (u[6]), .A (n_0_67), .B (y[6]));
XNOR2_X2 i_0_105 (.ZN (n_0_66), .A (z[5]), .B (x[5]));
XNOR2_X2 i_0_104 (.ZN (u[5]), .A (y[5]), .B (n_0_66));
XNOR2_X1 i_0_103 (.ZN (n_0_65), .A (z[4]), .B (x[4]));
XNOR2_X1 i_0_102 (.ZN (u[4]), .A (y[4]), .B (n_0_65));
XNOR2_X1 i_0_101 (.ZN (n_0_64), .A (z[3]), .B (x[3]));
XNOR2_X1 i_0_100 (.ZN (u[3]), .A (y[3]), .B (n_0_64));
XOR2_X1 i_0_99 (.Z (u[2]), .A (y[2]), .B (x[2]));
NOR2_X1 i_0_98 (.ZN (n_0_63), .A1 (y[61]), .A2 (x[61]));
NAND2_X1 i_0_97 (.ZN (n_0_62), .A1 (y[61]), .A2 (x[61]));
AOI21_X1 i_0_96 (.ZN (v[62]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_98));
AOI21_X1 i_0_95 (.ZN (v[36]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_97));
AOI21_X1 i_0_94 (.ZN (v[35]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_96));
NAND2_X1 i_0_93 (.ZN (n_0_61), .A1 (z[33]), .A2 (x[61]));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (y[33]), .B1 (z[33]), .B2 (x[61]));
NAND2_X1 i_0_91 (.ZN (v[34]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_88 (.ZN (v[33]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_85 (.ZN (v[32]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_82 (.ZN (v[31]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_79 (.ZN (v[30]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_76 (.ZN (v[29]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_73 (.ZN (v[28]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_70 (.ZN (v[27]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_67 (.ZN (v[26]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_64 (.ZN (v[25]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_61 (.ZN (v[24]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_58 (.ZN (v[23]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_55 (.ZN (v[22]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_52 (.ZN (v[21]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_49 (.ZN (v[20]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_46 (.ZN (v[19]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_43 (.ZN (v[18]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_40 (.ZN (v[17]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_37 (.ZN (v[16]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_34 (.ZN (v[15]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X2 i_0_31 (.ZN (v[14]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X4 i_0_28 (.ZN (v[13]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X2 i_0_25 (.ZN (v[12]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[10]), .A2 (x[10]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[10]), .B1 (z[10]), .B2 (x[10]));
NAND2_X1 i_0_22 (.ZN (v[11]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[9]), .A2 (x[9]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[9]), .B1 (z[9]), .B2 (x[9]));
NAND2_X1 i_0_19 (.ZN (v[10]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[8]), .A2 (x[8]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[8]), .B1 (z[8]), .B2 (x[8]));
NAND2_X1 i_0_16 (.ZN (v[9]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[7]), .A2 (x[7]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[7]), .B1 (z[7]), .B2 (x[7]));
NAND2_X1 i_0_13 (.ZN (v[8]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[6]), .A2 (x[6]));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[5]), .A2 (x[5]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[5]), .B1 (z[5]), .B2 (x[5]));
NAND2_X1 i_0_7 (.ZN (v[6]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[4]), .A2 (x[4]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[4]), .B1 (z[4]), .B2 (x[4]));
NAND2_X1 i_0_4 (.ZN (v[5]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[3]), .A2 (x[3]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[3]), .B1 (z[3]), .B2 (x[3]));
NAND2_X1 i_0_1 (.ZN (v[4]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[3]), .A1 (y[2]), .A2 (x[2]));
OAI21_X2 slo__mro_c1 (.ZN (slo__mro_n3), .A (y[6]), .B1 (x[6]), .B2 (z[6]));
NAND2_X2 slo__mro_c2 (.ZN (v[7]), .A1 (slo__mro_n3), .A2 (n_0_7));

endmodule //CSA__3_5

module CSA__3_2 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire drc_ipo_n3;
wire slo__mro_n6;


INV_X1 i_0_245 (.ZN (n_0_124), .A (z[62]));
INV_X1 i_0_244 (.ZN (n_0_123), .A (z[61]));
INV_X1 i_0_243 (.ZN (n_0_122), .A (z[60]));
INV_X1 i_0_242 (.ZN (n_0_121), .A (z[59]));
INV_X1 i_0_241 (.ZN (n_0_120), .A (z[58]));
INV_X1 i_0_240 (.ZN (n_0_119), .A (z[57]));
INV_X1 i_0_239 (.ZN (n_0_118), .A (z[56]));
INV_X1 i_0_238 (.ZN (n_0_117), .A (z[55]));
INV_X1 i_0_237 (.ZN (n_0_116), .A (z[54]));
INV_X1 i_0_236 (.ZN (n_0_115), .A (z[53]));
INV_X1 i_0_235 (.ZN (n_0_114), .A (z[52]));
INV_X1 i_0_234 (.ZN (n_0_113), .A (z[51]));
INV_X1 i_0_233 (.ZN (n_0_112), .A (z[50]));
INV_X1 i_0_232 (.ZN (n_0_111), .A (z[49]));
INV_X1 i_0_231 (.ZN (n_0_110), .A (z[48]));
INV_X1 i_0_230 (.ZN (n_0_109), .A (z[47]));
INV_X1 i_0_229 (.ZN (n_0_108), .A (z[46]));
INV_X1 i_0_228 (.ZN (n_0_107), .A (z[45]));
INV_X1 i_0_227 (.ZN (n_0_106), .A (z[44]));
INV_X1 i_0_226 (.ZN (n_0_105), .A (z[43]));
INV_X1 i_0_225 (.ZN (n_0_104), .A (z[42]));
INV_X1 i_0_224 (.ZN (n_0_103), .A (z[41]));
INV_X1 i_0_223 (.ZN (n_0_102), .A (z[40]));
INV_X1 i_0_222 (.ZN (n_0_101), .A (z[39]));
INV_X1 i_0_221 (.ZN (n_0_100), .A (z[38]));
INV_X1 i_0_220 (.ZN (n_0_99), .A (z[37]));
XOR2_X1 i_0_219 (.Z (n_0_98), .A (y[62]), .B (x[62]));
XOR2_X1 i_0_218 (.Z (u[63]), .A (z[63]), .B (drc_ipo_n3));
XNOR2_X1 i_0_217 (.ZN (u[62]), .A (n_0_124), .B (drc_ipo_n3));
XNOR2_X1 i_0_216 (.ZN (u[61]), .A (n_0_123), .B (drc_ipo_n3));
XNOR2_X1 i_0_215 (.ZN (u[60]), .A (n_0_122), .B (drc_ipo_n3));
XNOR2_X1 i_0_214 (.ZN (u[59]), .A (n_0_121), .B (drc_ipo_n3));
XNOR2_X1 i_0_213 (.ZN (u[58]), .A (n_0_120), .B (drc_ipo_n3));
XNOR2_X1 i_0_212 (.ZN (u[57]), .A (n_0_119), .B (drc_ipo_n3));
XNOR2_X1 i_0_211 (.ZN (u[56]), .A (n_0_118), .B (drc_ipo_n3));
XNOR2_X1 i_0_210 (.ZN (u[55]), .A (n_0_117), .B (drc_ipo_n3));
XNOR2_X1 i_0_209 (.ZN (u[54]), .A (n_0_116), .B (drc_ipo_n3));
XNOR2_X1 i_0_208 (.ZN (u[53]), .A (n_0_115), .B (drc_ipo_n3));
XNOR2_X1 i_0_207 (.ZN (u[52]), .A (n_0_114), .B (drc_ipo_n3));
XNOR2_X1 i_0_206 (.ZN (u[51]), .A (n_0_113), .B (drc_ipo_n3));
XNOR2_X1 i_0_205 (.ZN (u[50]), .A (n_0_112), .B (drc_ipo_n3));
XNOR2_X1 i_0_204 (.ZN (u[49]), .A (n_0_111), .B (drc_ipo_n3));
XNOR2_X1 i_0_203 (.ZN (u[48]), .A (n_0_110), .B (drc_ipo_n3));
XNOR2_X1 i_0_202 (.ZN (u[47]), .A (n_0_109), .B (drc_ipo_n3));
XNOR2_X1 i_0_201 (.ZN (u[46]), .A (n_0_108), .B (drc_ipo_n3));
XNOR2_X1 i_0_200 (.ZN (u[45]), .A (n_0_107), .B (drc_ipo_n3));
XNOR2_X1 i_0_199 (.ZN (u[44]), .A (n_0_106), .B (drc_ipo_n3));
XNOR2_X1 i_0_198 (.ZN (u[43]), .A (n_0_105), .B (drc_ipo_n3));
XNOR2_X1 i_0_197 (.ZN (u[42]), .A (n_0_104), .B (drc_ipo_n3));
XNOR2_X1 i_0_196 (.ZN (u[41]), .A (n_0_103), .B (drc_ipo_n3));
XNOR2_X1 i_0_195 (.ZN (u[40]), .A (n_0_102), .B (drc_ipo_n3));
XNOR2_X1 i_0_194 (.ZN (u[39]), .A (n_0_101), .B (drc_ipo_n3));
XNOR2_X1 i_0_193 (.ZN (u[38]), .A (n_0_100), .B (drc_ipo_n3));
XNOR2_X1 i_0_192 (.ZN (u[37]), .A (n_0_99), .B (drc_ipo_n3));
XNOR2_X1 i_0_191 (.ZN (n_0_97), .A (z[36]), .B (x[62]));
XNOR2_X2 i_0_190 (.ZN (u[36]), .A (y[36]), .B (n_0_97));
XNOR2_X1 i_0_189 (.ZN (n_0_96), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_188 (.ZN (u[35]), .A (y[35]), .B (n_0_96));
XNOR2_X1 i_0_187 (.ZN (n_0_95), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_186 (.ZN (u[34]), .A (y[34]), .B (n_0_95));
XNOR2_X1 i_0_185 (.ZN (n_0_94), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_184 (.ZN (u[33]), .A (y[33]), .B (n_0_94));
XNOR2_X1 i_0_183 (.ZN (n_0_93), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_182 (.ZN (u[32]), .A (y[32]), .B (n_0_93));
XNOR2_X1 i_0_181 (.ZN (n_0_92), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_180 (.ZN (u[31]), .A (y[31]), .B (n_0_92));
XNOR2_X1 i_0_179 (.ZN (n_0_91), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_178 (.ZN (u[30]), .A (y[30]), .B (n_0_91));
XNOR2_X1 i_0_177 (.ZN (n_0_90), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_176 (.ZN (u[29]), .A (y[29]), .B (n_0_90));
XNOR2_X1 i_0_175 (.ZN (n_0_89), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_174 (.ZN (u[28]), .A (y[28]), .B (n_0_89));
XNOR2_X1 i_0_173 (.ZN (n_0_88), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_172 (.ZN (u[27]), .A (y[27]), .B (n_0_88));
XNOR2_X1 i_0_171 (.ZN (n_0_87), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_170 (.ZN (u[26]), .A (y[26]), .B (n_0_87));
XNOR2_X1 i_0_169 (.ZN (n_0_86), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_168 (.ZN (u[25]), .A (y[25]), .B (n_0_86));
XNOR2_X1 i_0_167 (.ZN (n_0_85), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_166 (.ZN (u[24]), .A (y[24]), .B (n_0_85));
XNOR2_X1 i_0_165 (.ZN (n_0_84), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_164 (.ZN (u[23]), .A (y[23]), .B (n_0_84));
XNOR2_X1 i_0_163 (.ZN (n_0_83), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_162 (.ZN (u[22]), .A (y[22]), .B (n_0_83));
XNOR2_X1 i_0_161 (.ZN (n_0_82), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_160 (.ZN (u[21]), .A (y[21]), .B (n_0_82));
XNOR2_X1 i_0_159 (.ZN (n_0_81), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_158 (.ZN (u[20]), .A (y[20]), .B (n_0_81));
XNOR2_X1 i_0_157 (.ZN (n_0_80), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_156 (.ZN (u[19]), .A (y[19]), .B (n_0_80));
XNOR2_X1 i_0_155 (.ZN (n_0_79), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_154 (.ZN (u[18]), .A (y[18]), .B (n_0_79));
XNOR2_X1 i_0_153 (.ZN (n_0_78), .A (z[17]), .B (x[17]));
XNOR2_X2 i_0_152 (.ZN (u[17]), .A (y[17]), .B (n_0_78));
XNOR2_X1 i_0_151 (.ZN (n_0_77), .A (z[16]), .B (x[16]));
XNOR2_X2 i_0_150 (.ZN (u[16]), .A (y[16]), .B (n_0_77));
XNOR2_X2 i_0_149 (.ZN (n_0_76), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_148 (.ZN (u[15]), .A (y[15]), .B (n_0_76));
XNOR2_X2 i_0_147 (.ZN (n_0_75), .A (z[14]), .B (x[14]));
XNOR2_X2 i_0_146 (.ZN (u[14]), .A (y[14]), .B (n_0_75));
XNOR2_X2 i_0_145 (.ZN (n_0_74), .A (z[13]), .B (x[13]));
XNOR2_X2 i_0_144 (.ZN (u[13]), .A (n_0_74), .B (y[13]));
XNOR2_X2 i_0_143 (.ZN (n_0_73), .A (x[12]), .B (z[12]));
XNOR2_X2 i_0_142 (.ZN (u[12]), .A (n_0_73), .B (y[12]));
XNOR2_X2 i_0_141 (.ZN (n_0_72), .A (x[11]), .B (z[11]));
XNOR2_X2 i_0_140 (.ZN (u[11]), .A (n_0_72), .B (y[11]));
XNOR2_X2 i_0_139 (.ZN (n_0_71), .A (z[10]), .B (x[10]));
XNOR2_X2 i_0_138 (.ZN (u[10]), .A (n_0_71), .B (y[10]));
XNOR2_X2 i_0_135 (.ZN (n_0_69), .A (x[8]), .B (z[8]));
XNOR2_X2 i_0_134 (.ZN (u[8]), .A (n_0_69), .B (y[8]));
XNOR2_X2 i_0_133 (.ZN (n_0_68), .A (z[7]), .B (x[7]));
XNOR2_X2 i_0_132 (.ZN (u[7]), .A (n_0_68), .B (y[7]));
XNOR2_X2 i_0_131 (.ZN (n_0_67), .A (z[6]), .B (x[6]));
XNOR2_X2 i_0_130 (.ZN (u[6]), .A (y[6]), .B (n_0_67));
XNOR2_X2 i_0_129 (.ZN (n_0_66), .A (z[5]), .B (x[5]));
XNOR2_X2 i_0_128 (.ZN (u[5]), .A (y[5]), .B (n_0_66));
XOR2_X1 i_0_127 (.Z (u[4]), .A (y[4]), .B (x[4]));
XOR2_X1 i_0_126 (.Z (u[3]), .A (y[3]), .B (x[3]));
NAND2_X2 i_0_125 (.ZN (n_0_65), .A1 (y[62]), .A2 (x[62]));
NOR2_X4 i_0_124 (.ZN (n_0_64), .A1 (y[62]), .A2 (x[62]));
OAI21_X1 i_0_123 (.ZN (v[63]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_124));
OAI21_X1 i_0_122 (.ZN (v[62]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_123));
OAI21_X1 i_0_121 (.ZN (v[61]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_122));
OAI21_X1 i_0_120 (.ZN (v[60]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_121));
OAI21_X1 i_0_119 (.ZN (v[59]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_120));
OAI21_X1 i_0_118 (.ZN (v[58]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_119));
OAI21_X1 i_0_117 (.ZN (v[57]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_118));
OAI21_X1 i_0_116 (.ZN (v[56]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_117));
OAI21_X1 i_0_115 (.ZN (v[55]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_116));
OAI21_X1 i_0_114 (.ZN (v[54]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_115));
OAI21_X1 i_0_113 (.ZN (v[53]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_114));
OAI21_X1 i_0_112 (.ZN (v[52]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_113));
OAI21_X1 i_0_111 (.ZN (v[51]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_112));
OAI21_X1 i_0_110 (.ZN (v[50]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_111));
OAI21_X1 i_0_109 (.ZN (v[49]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_110));
OAI21_X1 i_0_108 (.ZN (v[48]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_109));
OAI21_X1 i_0_107 (.ZN (v[47]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_108));
OAI21_X1 i_0_106 (.ZN (v[46]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_107));
OAI21_X1 i_0_105 (.ZN (v[45]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_106));
OAI21_X1 i_0_104 (.ZN (v[44]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_105));
OAI21_X1 i_0_103 (.ZN (v[43]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_104));
OAI21_X1 i_0_102 (.ZN (v[42]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_103));
OAI21_X1 i_0_101 (.ZN (v[41]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_102));
OAI21_X1 i_0_100 (.ZN (v[40]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_101));
OAI21_X1 i_0_99 (.ZN (v[39]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_100));
OAI21_X1 i_0_98 (.ZN (v[38]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_99));
NAND2_X1 i_0_97 (.ZN (n_0_63), .A1 (z[36]), .A2 (x[62]));
OAI21_X1 i_0_96 (.ZN (n_0_62), .A (y[36]), .B1 (z[36]), .B2 (x[62]));
NAND2_X1 i_0_95 (.ZN (v[37]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_94 (.ZN (n_0_61), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_93 (.ZN (n_0_60), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_92 (.ZN (v[36]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_91 (.ZN (n_0_59), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_90 (.ZN (n_0_58), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_89 (.ZN (v[35]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_88 (.ZN (n_0_57), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_87 (.ZN (n_0_56), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_86 (.ZN (v[34]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_85 (.ZN (n_0_55), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_84 (.ZN (n_0_54), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_83 (.ZN (v[33]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_82 (.ZN (n_0_53), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_81 (.ZN (n_0_52), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_80 (.ZN (v[32]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_79 (.ZN (n_0_51), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_78 (.ZN (n_0_50), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_77 (.ZN (v[31]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_76 (.ZN (n_0_49), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_75 (.ZN (n_0_48), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_74 (.ZN (v[30]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_73 (.ZN (n_0_47), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_72 (.ZN (n_0_46), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_71 (.ZN (v[29]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_70 (.ZN (n_0_45), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_69 (.ZN (n_0_44), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_68 (.ZN (v[28]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_67 (.ZN (n_0_43), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_66 (.ZN (n_0_42), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_65 (.ZN (v[27]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_64 (.ZN (n_0_41), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_63 (.ZN (n_0_40), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_62 (.ZN (v[26]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_61 (.ZN (n_0_39), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_60 (.ZN (n_0_38), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_59 (.ZN (v[25]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_58 (.ZN (n_0_37), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_57 (.ZN (n_0_36), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_56 (.ZN (v[24]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_55 (.ZN (n_0_35), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_54 (.ZN (n_0_34), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_53 (.ZN (v[23]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_52 (.ZN (n_0_33), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_51 (.ZN (n_0_32), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_50 (.ZN (v[22]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_49 (.ZN (n_0_31), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_48 (.ZN (n_0_30), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_47 (.ZN (v[21]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_46 (.ZN (n_0_29), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_45 (.ZN (n_0_28), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_44 (.ZN (v[20]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_43 (.ZN (n_0_27), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_42 (.ZN (n_0_26), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_41 (.ZN (v[19]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_40 (.ZN (n_0_25), .A1 (y[17]), .A2 (z[17]));
OAI21_X1 i_0_39 (.ZN (n_0_24), .A (x[17]), .B1 (z[17]), .B2 (y[17]));
NAND2_X1 i_0_38 (.ZN (v[18]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_37 (.ZN (n_0_23), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_36 (.ZN (n_0_22), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_35 (.ZN (v[17]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_34 (.ZN (n_0_21), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_33 (.ZN (n_0_20), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_32 (.ZN (v[16]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_31 (.ZN (n_0_19), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_30 (.ZN (n_0_18), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_29 (.ZN (v[15]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_28 (.ZN (n_0_17), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_27 (.ZN (n_0_16), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X2 i_0_26 (.ZN (v[14]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_25 (.ZN (n_0_15), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_24 (.ZN (n_0_14), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X4 i_0_23 (.ZN (v[13]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_22 (.ZN (n_0_13), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_21 (.ZN (n_0_12), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X1 i_0_20 (.ZN (v[12]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_19 (.ZN (n_0_11), .A1 (z[10]), .A2 (x[10]));
OAI21_X1 i_0_18 (.ZN (n_0_10), .A (y[10]), .B1 (z[10]), .B2 (x[10]));
NAND2_X1 i_0_17 (.ZN (v[11]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_16 (.ZN (n_0_9), .A1 (z[9]), .A2 (x[9]));
OAI21_X1 i_0_15 (.ZN (n_0_8), .A (y[9]), .B1 (z[9]), .B2 (x[9]));
NAND2_X1 i_0_14 (.ZN (v[10]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_13 (.ZN (n_0_7), .A1 (z[8]), .A2 (x[8]));
OAI21_X1 i_0_12 (.ZN (n_0_6), .A (y[8]), .B1 (z[8]), .B2 (x[8]));
NAND2_X1 i_0_11 (.ZN (v[9]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_10 (.ZN (n_0_5), .A1 (z[7]), .A2 (x[7]));
OAI21_X1 i_0_9 (.ZN (n_0_4), .A (y[7]), .B1 (z[7]), .B2 (x[7]));
NAND2_X2 i_0_8 (.ZN (v[8]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_7 (.ZN (n_0_3), .A1 (z[6]), .A2 (x[6]));
OAI21_X1 i_0_6 (.ZN (n_0_2), .A (y[6]), .B1 (z[6]), .B2 (x[6]));
NAND2_X1 i_0_5 (.ZN (v[7]), .A1 (n_0_2), .A2 (n_0_3));
NAND2_X1 i_0_4 (.ZN (n_0_1), .A1 (z[5]), .A2 (x[5]));
OAI21_X1 i_0_3 (.ZN (n_0_0), .A (y[5]), .B1 (z[5]), .B2 (x[5]));
NAND2_X2 i_0_2 (.ZN (v[6]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X2 i_0_1 (.ZN (v[5]), .A1 (y[4]), .A2 (x[4]));
AND2_X1 i_0_0 (.ZN (v[4]), .A1 (y[3]), .A2 (x[3]));
CLKBUF_X3 drc_ipo_c3 (.Z (drc_ipo_n3), .A (n_0_98));
XNOR2_X2 slo__mro_c4 (.ZN (slo__mro_n6), .A (z[9]), .B (y[9]));
XNOR2_X2 slo__mro_c5 (.ZN (u[9]), .A (slo__mro_n6), .B (x[9]));

endmodule //CSA__3_2

module CSA__0_72 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire drc_ipo_n3;


INV_X1 i_0_230 (.ZN (n_0_121), .A (x[62]));
INV_X1 i_0_229 (.ZN (n_0_120), .A (x[61]));
INV_X1 i_0_228 (.ZN (n_0_119), .A (x[60]));
INV_X1 i_0_227 (.ZN (n_0_118), .A (x[59]));
INV_X1 i_0_226 (.ZN (n_0_117), .A (x[58]));
INV_X1 i_0_225 (.ZN (n_0_116), .A (x[57]));
INV_X1 i_0_224 (.ZN (n_0_115), .A (x[56]));
INV_X1 i_0_223 (.ZN (n_0_114), .A (x[55]));
INV_X1 i_0_222 (.ZN (n_0_113), .A (x[54]));
INV_X1 i_0_221 (.ZN (n_0_112), .A (x[53]));
INV_X1 i_0_220 (.ZN (n_0_111), .A (x[52]));
INV_X1 i_0_219 (.ZN (n_0_110), .A (x[51]));
INV_X1 i_0_218 (.ZN (n_0_109), .A (x[50]));
INV_X1 i_0_217 (.ZN (n_0_108), .A (x[49]));
INV_X1 i_0_216 (.ZN (n_0_107), .A (x[48]));
INV_X1 i_0_215 (.ZN (n_0_106), .A (x[47]));
INV_X1 i_0_214 (.ZN (n_0_105), .A (x[46]));
XOR2_X1 i_0_213 (.Z (n_0_104), .A (y[63]), .B (z[63]));
XOR2_X1 i_0_212 (.Z (u[63]), .A (x[63]), .B (drc_ipo_n3));
XNOR2_X1 i_0_211 (.ZN (u[62]), .A (n_0_121), .B (drc_ipo_n3));
XNOR2_X1 i_0_210 (.ZN (u[61]), .A (n_0_120), .B (drc_ipo_n3));
XNOR2_X1 i_0_209 (.ZN (u[60]), .A (n_0_119), .B (drc_ipo_n3));
XNOR2_X1 i_0_208 (.ZN (u[59]), .A (n_0_118), .B (drc_ipo_n3));
XNOR2_X1 i_0_207 (.ZN (u[58]), .A (n_0_117), .B (drc_ipo_n3));
XNOR2_X1 i_0_206 (.ZN (u[57]), .A (n_0_116), .B (drc_ipo_n3));
XNOR2_X1 i_0_205 (.ZN (u[56]), .A (n_0_115), .B (drc_ipo_n3));
XNOR2_X1 i_0_204 (.ZN (u[55]), .A (n_0_114), .B (drc_ipo_n3));
XNOR2_X1 i_0_203 (.ZN (u[54]), .A (n_0_113), .B (drc_ipo_n3));
XNOR2_X1 i_0_202 (.ZN (u[53]), .A (n_0_112), .B (drc_ipo_n3));
XNOR2_X1 i_0_201 (.ZN (u[52]), .A (n_0_111), .B (drc_ipo_n3));
XNOR2_X1 i_0_200 (.ZN (u[51]), .A (n_0_110), .B (drc_ipo_n3));
XNOR2_X1 i_0_199 (.ZN (u[50]), .A (n_0_109), .B (drc_ipo_n3));
XNOR2_X1 i_0_198 (.ZN (u[49]), .A (n_0_108), .B (drc_ipo_n3));
XNOR2_X1 i_0_197 (.ZN (u[48]), .A (n_0_107), .B (drc_ipo_n3));
XNOR2_X1 i_0_196 (.ZN (u[47]), .A (n_0_106), .B (drc_ipo_n3));
XNOR2_X1 i_0_195 (.ZN (u[46]), .A (n_0_105), .B (drc_ipo_n3));
XNOR2_X1 i_0_194 (.ZN (n_0_103), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_193 (.ZN (u[45]), .A (y[63]), .B (n_0_103));
XNOR2_X1 i_0_192 (.ZN (n_0_102), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_191 (.ZN (u[44]), .A (y[44]), .B (n_0_102));
XNOR2_X1 i_0_190 (.ZN (n_0_101), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_189 (.ZN (u[43]), .A (y[43]), .B (n_0_101));
XNOR2_X1 i_0_188 (.ZN (n_0_100), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_187 (.ZN (u[42]), .A (y[42]), .B (n_0_100));
XNOR2_X1 i_0_186 (.ZN (n_0_99), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_185 (.ZN (u[41]), .A (y[41]), .B (n_0_99));
XNOR2_X1 i_0_184 (.ZN (n_0_98), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_183 (.ZN (u[40]), .A (y[40]), .B (n_0_98));
XNOR2_X1 i_0_182 (.ZN (n_0_97), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_181 (.ZN (u[39]), .A (y[39]), .B (n_0_97));
XNOR2_X1 i_0_180 (.ZN (n_0_96), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_179 (.ZN (u[38]), .A (y[38]), .B (n_0_96));
XNOR2_X1 i_0_178 (.ZN (n_0_95), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_177 (.ZN (u[37]), .A (y[37]), .B (n_0_95));
XNOR2_X1 i_0_176 (.ZN (n_0_94), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_175 (.ZN (u[36]), .A (y[36]), .B (n_0_94));
XNOR2_X1 i_0_174 (.ZN (n_0_93), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_173 (.ZN (u[35]), .A (y[35]), .B (n_0_93));
XNOR2_X1 i_0_172 (.ZN (n_0_92), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_171 (.ZN (u[34]), .A (y[34]), .B (n_0_92));
XNOR2_X1 i_0_170 (.ZN (n_0_91), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_169 (.ZN (u[33]), .A (y[33]), .B (n_0_91));
XNOR2_X1 i_0_168 (.ZN (n_0_90), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_167 (.ZN (u[32]), .A (y[32]), .B (n_0_90));
XNOR2_X1 i_0_166 (.ZN (n_0_89), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_165 (.ZN (u[31]), .A (y[31]), .B (n_0_89));
XNOR2_X1 i_0_164 (.ZN (n_0_88), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_163 (.ZN (u[30]), .A (y[30]), .B (n_0_88));
XNOR2_X1 i_0_162 (.ZN (n_0_87), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_161 (.ZN (u[29]), .A (y[29]), .B (n_0_87));
XNOR2_X1 i_0_160 (.ZN (n_0_86), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_159 (.ZN (u[28]), .A (y[28]), .B (n_0_86));
XNOR2_X1 i_0_158 (.ZN (n_0_85), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_157 (.ZN (u[27]), .A (y[27]), .B (n_0_85));
XNOR2_X1 i_0_156 (.ZN (n_0_84), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_155 (.ZN (u[26]), .A (y[26]), .B (n_0_84));
XNOR2_X1 i_0_154 (.ZN (n_0_83), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_153 (.ZN (u[25]), .A (y[25]), .B (n_0_83));
XNOR2_X1 i_0_152 (.ZN (n_0_82), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_151 (.ZN (u[24]), .A (y[24]), .B (n_0_82));
XNOR2_X1 i_0_150 (.ZN (n_0_81), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_149 (.ZN (u[23]), .A (y[23]), .B (n_0_81));
XNOR2_X1 i_0_148 (.ZN (n_0_80), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_147 (.ZN (u[22]), .A (y[22]), .B (n_0_80));
XNOR2_X1 i_0_146 (.ZN (n_0_79), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_145 (.ZN (u[21]), .A (y[21]), .B (n_0_79));
XNOR2_X1 i_0_144 (.ZN (n_0_78), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_143 (.ZN (u[20]), .A (y[20]), .B (n_0_78));
XNOR2_X1 i_0_142 (.ZN (n_0_77), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_141 (.ZN (u[19]), .A (y[19]), .B (n_0_77));
XNOR2_X1 i_0_140 (.ZN (n_0_76), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_139 (.ZN (u[18]), .A (y[18]), .B (n_0_76));
XNOR2_X1 i_0_138 (.ZN (n_0_75), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_137 (.ZN (u[17]), .A (y[17]), .B (n_0_75));
XNOR2_X1 i_0_136 (.ZN (n_0_74), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_135 (.ZN (u[16]), .A (y[16]), .B (n_0_74));
XNOR2_X2 i_0_134 (.ZN (n_0_73), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_133 (.ZN (u[15]), .A (y[15]), .B (n_0_73));
XNOR2_X2 i_0_132 (.ZN (n_0_72), .A (z[14]), .B (x[14]));
XNOR2_X2 i_0_131 (.ZN (u[14]), .A (y[14]), .B (n_0_72));
XNOR2_X1 i_0_130 (.ZN (n_0_71), .A (z[13]), .B (x[13]));
XNOR2_X2 i_0_129 (.ZN (u[13]), .A (y[13]), .B (n_0_71));
XNOR2_X1 i_0_128 (.ZN (n_0_70), .A (z[12]), .B (x[12]));
XNOR2_X2 i_0_127 (.ZN (u[12]), .A (y[12]), .B (n_0_70));
XOR2_X2 i_0_126 (.Z (u[11]), .A (y[11]), .B (x[11]));
XOR2_X2 i_0_125 (.Z (u[10]), .A (y[10]), .B (x[10]));
XOR2_X1 i_0_124 (.Z (u[9]), .A (y[9]), .B (x[9]));
NAND2_X1 i_0_123 (.ZN (n_0_69), .A1 (y[63]), .A2 (z[63]));
NOR2_X2 i_0_122 (.ZN (n_0_68), .A1 (y[63]), .A2 (z[63]));
OAI21_X1 i_0_121 (.ZN (v[63]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_121));
OAI21_X1 i_0_120 (.ZN (v[62]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_120));
OAI21_X1 i_0_119 (.ZN (v[61]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_119));
OAI21_X1 i_0_118 (.ZN (v[60]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_118));
OAI21_X1 i_0_117 (.ZN (v[59]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_117));
OAI21_X1 i_0_116 (.ZN (v[58]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_116));
OAI21_X1 i_0_115 (.ZN (v[57]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_115));
OAI21_X1 i_0_114 (.ZN (v[56]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_114));
OAI21_X1 i_0_113 (.ZN (v[55]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_113));
OAI21_X1 i_0_112 (.ZN (v[54]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_112));
OAI21_X1 i_0_111 (.ZN (v[53]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_111));
OAI21_X1 i_0_110 (.ZN (v[52]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_110));
OAI21_X1 i_0_109 (.ZN (v[51]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_109));
OAI21_X1 i_0_108 (.ZN (v[50]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_108));
OAI21_X1 i_0_107 (.ZN (v[49]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_107));
OAI21_X1 i_0_106 (.ZN (v[48]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_106));
OAI21_X1 i_0_105 (.ZN (v[47]), .A (n_0_69), .B1 (n_0_68), .B2 (n_0_105));
NAND2_X1 i_0_104 (.ZN (n_0_67), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_103 (.ZN (n_0_66), .A (y[63]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_102 (.ZN (v[46]), .A1 (n_0_67), .A2 (n_0_66));
NAND2_X1 i_0_101 (.ZN (n_0_65), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_100 (.ZN (n_0_64), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_99 (.ZN (v[45]), .A1 (n_0_65), .A2 (n_0_64));
NAND2_X1 i_0_98 (.ZN (n_0_63), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_97 (.ZN (n_0_62), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_96 (.ZN (v[44]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_95 (.ZN (n_0_61), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_94 (.ZN (n_0_60), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_93 (.ZN (v[43]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_92 (.ZN (n_0_59), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_91 (.ZN (n_0_58), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_90 (.ZN (v[42]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_89 (.ZN (n_0_57), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_88 (.ZN (n_0_56), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_87 (.ZN (v[41]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_86 (.ZN (n_0_55), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_85 (.ZN (n_0_54), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_84 (.ZN (v[40]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_83 (.ZN (n_0_53), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_82 (.ZN (n_0_52), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_81 (.ZN (v[39]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_80 (.ZN (n_0_51), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_79 (.ZN (n_0_50), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_78 (.ZN (v[38]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_77 (.ZN (n_0_49), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_76 (.ZN (n_0_48), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_75 (.ZN (v[37]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_74 (.ZN (n_0_47), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_73 (.ZN (n_0_46), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_72 (.ZN (v[36]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_71 (.ZN (n_0_45), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_70 (.ZN (n_0_44), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_69 (.ZN (v[35]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_68 (.ZN (n_0_43), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_67 (.ZN (n_0_42), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_66 (.ZN (v[34]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_65 (.ZN (n_0_41), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_64 (.ZN (n_0_40), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_63 (.ZN (v[33]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_62 (.ZN (n_0_39), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_61 (.ZN (n_0_38), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_60 (.ZN (v[32]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_59 (.ZN (n_0_37), .A1 (y[30]), .A2 (x[30]));
OAI21_X1 i_0_58 (.ZN (n_0_36), .A (z[30]), .B1 (x[30]), .B2 (y[30]));
NAND2_X1 i_0_57 (.ZN (v[31]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_56 (.ZN (n_0_35), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_55 (.ZN (n_0_34), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_54 (.ZN (v[30]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_53 (.ZN (n_0_33), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_52 (.ZN (n_0_32), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_51 (.ZN (v[29]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_50 (.ZN (n_0_31), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_49 (.ZN (n_0_30), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_48 (.ZN (v[28]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_47 (.ZN (n_0_29), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_46 (.ZN (n_0_28), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_45 (.ZN (v[27]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_44 (.ZN (n_0_27), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_43 (.ZN (n_0_26), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_42 (.ZN (v[26]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_41 (.ZN (n_0_25), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_40 (.ZN (n_0_24), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_39 (.ZN (v[25]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_38 (.ZN (n_0_23), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_37 (.ZN (n_0_22), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_36 (.ZN (v[24]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_35 (.ZN (n_0_21), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_34 (.ZN (n_0_20), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_33 (.ZN (v[23]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_32 (.ZN (n_0_19), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_31 (.ZN (n_0_18), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_30 (.ZN (v[22]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_29 (.ZN (n_0_17), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_28 (.ZN (n_0_16), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_27 (.ZN (v[21]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_26 (.ZN (n_0_15), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_25 (.ZN (n_0_14), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_24 (.ZN (v[20]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_23 (.ZN (n_0_13), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_22 (.ZN (n_0_12), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_21 (.ZN (v[19]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_20 (.ZN (n_0_11), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_19 (.ZN (n_0_10), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_18 (.ZN (v[18]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_17 (.ZN (n_0_9), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_16 (.ZN (n_0_8), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_15 (.ZN (v[17]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_14 (.ZN (n_0_7), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_13 (.ZN (n_0_6), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X2 i_0_12 (.ZN (v[16]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_11 (.ZN (n_0_5), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_10 (.ZN (n_0_4), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X4 i_0_9 (.ZN (v[15]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_8 (.ZN (n_0_3), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_7 (.ZN (n_0_2), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X1 i_0_6 (.ZN (v[14]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_5 (.ZN (n_0_1), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_4 (.ZN (n_0_0), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X1 i_0_3 (.ZN (v[13]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X2 i_0_2 (.ZN (v[12]), .A1 (y[11]), .A2 (x[11]));
AND2_X1 i_0_1 (.ZN (v[11]), .A1 (y[10]), .A2 (x[10]));
AND2_X1 i_0_0 (.ZN (v[10]), .A1 (y[9]), .A2 (x[9]));
BUF_X1 drc_ipo_c3 (.Z (drc_ipo_n3), .A (n_0_104));

endmodule //CSA__0_72

module CSA__2_11 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;


XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[62]), .B (x[62]));
XOR2_X1 i_0_158 (.Z (u[63]), .A (z[62]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[41]), .A (z[41]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[40]), .B (x[62]));
XNOR2_X1 i_0_155 (.ZN (u[40]), .A (y[40]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_153 (.ZN (u[39]), .A (y[39]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_151 (.ZN (u[38]), .A (y[38]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_149 (.ZN (u[37]), .A (y[37]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_147 (.ZN (u[36]), .A (y[36]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_145 (.ZN (u[35]), .A (y[35]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_143 (.ZN (u[34]), .A (y[34]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_141 (.ZN (u[33]), .A (y[33]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_139 (.ZN (u[32]), .A (y[32]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_137 (.ZN (u[31]), .A (y[31]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_135 (.ZN (u[30]), .A (y[30]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_133 (.ZN (u[29]), .A (y[29]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_131 (.ZN (u[28]), .A (y[28]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_129 (.ZN (u[27]), .A (y[27]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_127 (.ZN (u[26]), .A (y[26]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_125 (.ZN (u[25]), .A (y[25]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_123 (.ZN (u[24]), .A (y[24]), .B (n_0_76));
XNOR2_X1 i_0_122 (.ZN (n_0_75), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_121 (.ZN (u[23]), .A (y[23]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_119 (.ZN (u[22]), .A (y[22]), .B (n_0_74));
XNOR2_X1 i_0_118 (.ZN (n_0_73), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_117 (.ZN (u[21]), .A (y[21]), .B (n_0_73));
XNOR2_X1 i_0_116 (.ZN (n_0_72), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_115 (.ZN (u[20]), .A (y[20]), .B (n_0_72));
XNOR2_X1 i_0_114 (.ZN (n_0_71), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_113 (.ZN (u[19]), .A (y[19]), .B (n_0_71));
XNOR2_X1 i_0_112 (.ZN (n_0_70), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_111 (.ZN (u[18]), .A (y[18]), .B (n_0_70));
XNOR2_X1 i_0_110 (.ZN (n_0_69), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_109 (.ZN (u[17]), .A (y[17]), .B (n_0_69));
XNOR2_X1 i_0_108 (.ZN (n_0_68), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_107 (.ZN (u[16]), .A (y[16]), .B (n_0_68));
XNOR2_X2 i_0_106 (.ZN (n_0_67), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_105 (.ZN (u[15]), .A (y[15]), .B (n_0_67));
XNOR2_X1 i_0_104 (.ZN (n_0_66), .A (z[14]), .B (x[14]));
XNOR2_X1 i_0_103 (.ZN (u[14]), .A (y[14]), .B (n_0_66));
XNOR2_X2 i_0_102 (.ZN (n_0_65), .A (z[13]), .B (x[13]));
XNOR2_X1 i_0_101 (.ZN (u[13]), .A (y[13]), .B (n_0_65));
XNOR2_X2 i_0_100 (.ZN (n_0_64), .A (z[12]), .B (x[12]));
XNOR2_X2 i_0_99 (.ZN (u[12]), .A (n_0_64), .B (y[12]));
XNOR2_X2 i_0_98 (.ZN (n_0_63), .A (z[11]), .B (x[11]));
XNOR2_X2 i_0_97 (.ZN (u[11]), .A (n_0_63), .B (y[11]));
XOR2_X1 i_0_96 (.Z (u[10]), .A (y[10]), .B (x[10]));
NAND2_X1 i_0_95 (.ZN (n_0_62), .A1 (y[62]), .A2 (x[62]));
OAI21_X1 i_0_94 (.ZN (n_0_61), .A (z[62]), .B1 (x[62]), .B2 (y[62]));
NAND2_X1 i_0_93 (.ZN (v[63]), .A1 (n_0_62), .A2 (n_0_61));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (z[41]), .B1 (x[62]), .B2 (y[62]));
NAND2_X1 i_0_91 (.ZN (v[42]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[40]), .A2 (x[62]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[40]), .B1 (z[40]), .B2 (x[62]));
NAND2_X1 i_0_88 (.ZN (v[41]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_85 (.ZN (v[40]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_82 (.ZN (v[39]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_79 (.ZN (v[38]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_76 (.ZN (v[37]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_73 (.ZN (v[36]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_70 (.ZN (v[35]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_67 (.ZN (v[34]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_64 (.ZN (v[33]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_61 (.ZN (v[32]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_58 (.ZN (v[31]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_55 (.ZN (v[30]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_52 (.ZN (v[29]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_49 (.ZN (v[28]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_46 (.ZN (v[27]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_43 (.ZN (v[26]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_40 (.ZN (v[25]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_37 (.ZN (v[24]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_34 (.ZN (v[23]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_31 (.ZN (v[22]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_28 (.ZN (v[21]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_25 (.ZN (v[20]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_22 (.ZN (v[19]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_19 (.ZN (v[18]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_16 (.ZN (v[17]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_13 (.ZN (v[16]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_10 (.ZN (v[15]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X1 i_0_7 (.ZN (v[14]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X1 i_0_4 (.ZN (v[13]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X1 i_0_1 (.ZN (v[12]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[11]), .A1 (y[10]), .A2 (x[10]));

endmodule //CSA__2_11

module CSA__2_8 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire slo__sro_n3;


INV_X1 i_0_168 (.ZN (n_0_98), .A (z[63]));
INV_X1 i_0_167 (.ZN (n_0_97), .A (z[44]));
INV_X1 i_0_166 (.ZN (n_0_96), .A (z[43]));
XOR2_X1 i_0_165 (.Z (n_0_95), .A (y[63]), .B (x[63]));
XNOR2_X1 i_0_164 (.ZN (u[63]), .A (n_0_98), .B (n_0_95));
XNOR2_X1 i_0_163 (.ZN (u[44]), .A (n_0_97), .B (n_0_95));
XNOR2_X1 i_0_162 (.ZN (u[43]), .A (n_0_96), .B (n_0_95));
XNOR2_X1 i_0_161 (.ZN (n_0_94), .A (z[42]), .B (x[63]));
XNOR2_X1 i_0_160 (.ZN (u[42]), .A (y[42]), .B (n_0_94));
XNOR2_X1 i_0_159 (.ZN (n_0_93), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_158 (.ZN (u[41]), .A (y[41]), .B (n_0_93));
XNOR2_X1 i_0_157 (.ZN (n_0_92), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_156 (.ZN (u[40]), .A (y[40]), .B (n_0_92));
XNOR2_X1 i_0_155 (.ZN (n_0_91), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_154 (.ZN (u[39]), .A (y[39]), .B (n_0_91));
XNOR2_X1 i_0_153 (.ZN (n_0_90), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_152 (.ZN (u[38]), .A (y[38]), .B (n_0_90));
XNOR2_X1 i_0_151 (.ZN (n_0_89), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_150 (.ZN (u[37]), .A (y[37]), .B (n_0_89));
XNOR2_X1 i_0_149 (.ZN (n_0_88), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_148 (.ZN (u[36]), .A (y[36]), .B (n_0_88));
XNOR2_X1 i_0_147 (.ZN (n_0_87), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_146 (.ZN (u[35]), .A (y[35]), .B (n_0_87));
XNOR2_X1 i_0_145 (.ZN (n_0_86), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_144 (.ZN (u[34]), .A (y[34]), .B (n_0_86));
XNOR2_X1 i_0_143 (.ZN (n_0_85), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_142 (.ZN (u[33]), .A (y[33]), .B (n_0_85));
XNOR2_X1 i_0_141 (.ZN (n_0_84), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_140 (.ZN (u[32]), .A (y[32]), .B (n_0_84));
XNOR2_X1 i_0_139 (.ZN (n_0_83), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_138 (.ZN (u[31]), .A (y[31]), .B (n_0_83));
XNOR2_X1 i_0_137 (.ZN (n_0_82), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_136 (.ZN (u[30]), .A (y[30]), .B (n_0_82));
XNOR2_X1 i_0_135 (.ZN (n_0_81), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_134 (.ZN (u[29]), .A (y[29]), .B (n_0_81));
XNOR2_X1 i_0_133 (.ZN (n_0_80), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_132 (.ZN (u[28]), .A (y[28]), .B (n_0_80));
XNOR2_X1 i_0_131 (.ZN (n_0_79), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_130 (.ZN (u[27]), .A (y[27]), .B (n_0_79));
XNOR2_X1 i_0_129 (.ZN (n_0_78), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_128 (.ZN (u[26]), .A (y[26]), .B (n_0_78));
XNOR2_X1 i_0_127 (.ZN (n_0_77), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_126 (.ZN (u[25]), .A (y[25]), .B (n_0_77));
XNOR2_X1 i_0_125 (.ZN (n_0_76), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_124 (.ZN (u[24]), .A (y[24]), .B (n_0_76));
XNOR2_X1 i_0_123 (.ZN (n_0_75), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_122 (.ZN (u[23]), .A (y[23]), .B (n_0_75));
XNOR2_X1 i_0_121 (.ZN (n_0_74), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_120 (.ZN (u[22]), .A (y[22]), .B (n_0_74));
XNOR2_X1 i_0_119 (.ZN (n_0_73), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_118 (.ZN (u[21]), .A (y[21]), .B (n_0_73));
XNOR2_X1 i_0_117 (.ZN (n_0_72), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_116 (.ZN (u[20]), .A (y[20]), .B (n_0_72));
XNOR2_X1 i_0_115 (.ZN (n_0_71), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_114 (.ZN (u[19]), .A (y[19]), .B (n_0_71));
XNOR2_X1 i_0_113 (.ZN (n_0_70), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_112 (.ZN (u[18]), .A (y[18]), .B (n_0_70));
XNOR2_X1 i_0_111 (.ZN (n_0_69), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_110 (.ZN (u[17]), .A (y[17]), .B (n_0_69));
XNOR2_X1 i_0_109 (.ZN (n_0_68), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_108 (.ZN (u[16]), .A (y[16]), .B (n_0_68));
XNOR2_X1 i_0_107 (.ZN (n_0_67), .A (z[15]), .B (x[15]));
XNOR2_X1 i_0_106 (.ZN (u[15]), .A (y[15]), .B (n_0_67));
XNOR2_X2 i_0_105 (.ZN (n_0_66), .A (z[14]), .B (x[14]));
XNOR2_X2 i_0_104 (.ZN (u[14]), .A (y[14]), .B (n_0_66));
XNOR2_X2 i_0_103 (.ZN (n_0_65), .A (z[13]), .B (x[13]));
XNOR2_X1 i_0_102 (.ZN (u[13]), .A (y[13]), .B (n_0_65));
XNOR2_X2 i_0_101 (.ZN (n_0_64), .A (x[12]), .B (z[12]));
XNOR2_X2 i_0_100 (.ZN (u[12]), .A (n_0_64), .B (y[12]));
NOR2_X1 i_0_98 (.ZN (n_0_63), .A1 (y[63]), .A2 (x[63]));
NAND2_X1 i_0_97 (.ZN (n_0_62), .A1 (y[63]), .A2 (x[63]));
AOI21_X1 i_0_96 (.ZN (v[63]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_98));
AOI21_X1 i_0_95 (.ZN (v[45]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_97));
AOI21_X1 i_0_94 (.ZN (v[44]), .A (n_0_63), .B1 (n_0_62), .B2 (n_0_96));
NAND2_X1 i_0_93 (.ZN (n_0_61), .A1 (z[42]), .A2 (x[63]));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (y[42]), .B1 (z[42]), .B2 (x[63]));
NAND2_X1 i_0_91 (.ZN (v[43]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_88 (.ZN (v[42]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_85 (.ZN (v[41]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_82 (.ZN (v[40]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_79 (.ZN (v[39]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_76 (.ZN (v[38]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_73 (.ZN (v[37]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_70 (.ZN (v[36]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_67 (.ZN (v[35]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_64 (.ZN (v[34]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_61 (.ZN (v[33]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_58 (.ZN (v[32]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_55 (.ZN (v[31]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_52 (.ZN (v[30]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_49 (.ZN (v[29]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_46 (.ZN (v[28]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_43 (.ZN (v[27]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_40 (.ZN (v[26]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_37 (.ZN (v[25]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_34 (.ZN (v[24]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_31 (.ZN (v[23]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_28 (.ZN (v[22]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_25 (.ZN (v[21]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_22 (.ZN (v[20]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_19 (.ZN (v[19]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_16 (.ZN (v[18]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_13 (.ZN (v[17]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_10 (.ZN (v[16]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_7 (.ZN (v[15]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X1 i_0_4 (.ZN (v[14]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X1 i_0_1 (.ZN (v[13]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[12]), .A1 (y[11]), .A2 (x[11]));
INV_X1 slo__sro_c1 (.ZN (slo__sro_n3), .A (y[11]));
XNOR2_X1 slo__sro_c2 (.ZN (u[11]), .A (x[11]), .B (slo__sro_n3));

endmodule //CSA__2_8

module CSA__2_5 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire drc_ipo_n3;
wire slo__mro_n6;


INV_X1 i_0_236 (.ZN (n_0_121), .A (x[62]));
INV_X1 i_0_235 (.ZN (n_0_120), .A (x[61]));
INV_X1 i_0_234 (.ZN (n_0_119), .A (x[60]));
INV_X1 i_0_233 (.ZN (n_0_118), .A (x[59]));
INV_X1 i_0_232 (.ZN (n_0_117), .A (x[58]));
INV_X1 i_0_231 (.ZN (n_0_116), .A (x[57]));
INV_X1 i_0_230 (.ZN (n_0_115), .A (x[56]));
INV_X1 i_0_229 (.ZN (n_0_114), .A (x[55]));
INV_X1 i_0_228 (.ZN (n_0_113), .A (x[54]));
INV_X1 i_0_227 (.ZN (n_0_112), .A (x[53]));
INV_X1 i_0_226 (.ZN (n_0_111), .A (x[52]));
INV_X1 i_0_225 (.ZN (n_0_110), .A (x[51]));
INV_X1 i_0_224 (.ZN (n_0_109), .A (x[50]));
INV_X1 i_0_223 (.ZN (n_0_108), .A (x[49]));
INV_X1 i_0_222 (.ZN (n_0_107), .A (x[48]));
INV_X1 i_0_221 (.ZN (n_0_106), .A (x[47]));
INV_X1 i_0_220 (.ZN (n_0_105), .A (x[46]));
INV_X1 i_0_219 (.ZN (n_0_104), .A (x[45]));
INV_X1 i_0_218 (.ZN (n_0_103), .A (x[44]));
INV_X1 i_0_217 (.ZN (n_0_102), .A (x[43]));
INV_X1 i_0_216 (.ZN (n_0_101), .A (x[42]));
INV_X1 i_0_215 (.ZN (n_0_100), .A (x[41]));
INV_X1 i_0_214 (.ZN (n_0_99), .A (x[40]));
XOR2_X1 i_0_213 (.Z (n_0_98), .A (y[63]), .B (z[63]));
XOR2_X1 i_0_212 (.Z (u[63]), .A (x[63]), .B (drc_ipo_n3));
XNOR2_X1 i_0_211 (.ZN (u[62]), .A (n_0_121), .B (drc_ipo_n3));
XNOR2_X1 i_0_210 (.ZN (u[61]), .A (n_0_120), .B (drc_ipo_n3));
XNOR2_X1 i_0_209 (.ZN (u[60]), .A (n_0_119), .B (drc_ipo_n3));
XNOR2_X1 i_0_208 (.ZN (u[59]), .A (n_0_118), .B (drc_ipo_n3));
XNOR2_X1 i_0_207 (.ZN (u[58]), .A (n_0_117), .B (drc_ipo_n3));
XNOR2_X1 i_0_206 (.ZN (u[57]), .A (n_0_116), .B (drc_ipo_n3));
XNOR2_X1 i_0_205 (.ZN (u[56]), .A (n_0_115), .B (drc_ipo_n3));
XNOR2_X1 i_0_204 (.ZN (u[55]), .A (n_0_114), .B (drc_ipo_n3));
XNOR2_X1 i_0_203 (.ZN (u[54]), .A (n_0_113), .B (drc_ipo_n3));
XNOR2_X1 i_0_202 (.ZN (u[53]), .A (n_0_112), .B (drc_ipo_n3));
XNOR2_X1 i_0_201 (.ZN (u[52]), .A (n_0_111), .B (drc_ipo_n3));
XNOR2_X1 i_0_200 (.ZN (u[51]), .A (n_0_110), .B (drc_ipo_n3));
XNOR2_X1 i_0_199 (.ZN (u[50]), .A (n_0_109), .B (drc_ipo_n3));
XNOR2_X1 i_0_198 (.ZN (u[49]), .A (n_0_108), .B (drc_ipo_n3));
XNOR2_X1 i_0_197 (.ZN (u[48]), .A (n_0_107), .B (drc_ipo_n3));
XNOR2_X1 i_0_196 (.ZN (u[47]), .A (n_0_106), .B (drc_ipo_n3));
XNOR2_X1 i_0_195 (.ZN (u[46]), .A (n_0_105), .B (drc_ipo_n3));
XNOR2_X1 i_0_194 (.ZN (u[45]), .A (n_0_104), .B (drc_ipo_n3));
XNOR2_X1 i_0_193 (.ZN (u[44]), .A (n_0_103), .B (drc_ipo_n3));
XNOR2_X1 i_0_192 (.ZN (u[43]), .A (n_0_102), .B (drc_ipo_n3));
XNOR2_X1 i_0_191 (.ZN (u[42]), .A (n_0_101), .B (drc_ipo_n3));
XNOR2_X1 i_0_190 (.ZN (u[41]), .A (n_0_100), .B (drc_ipo_n3));
XNOR2_X1 i_0_189 (.ZN (u[40]), .A (n_0_99), .B (drc_ipo_n3));
XNOR2_X1 i_0_188 (.ZN (n_0_97), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_187 (.ZN (u[39]), .A (y[63]), .B (n_0_97));
XNOR2_X1 i_0_186 (.ZN (n_0_96), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_185 (.ZN (u[38]), .A (y[38]), .B (n_0_96));
XNOR2_X1 i_0_184 (.ZN (n_0_95), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_183 (.ZN (u[37]), .A (y[37]), .B (n_0_95));
XNOR2_X1 i_0_182 (.ZN (n_0_94), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_181 (.ZN (u[36]), .A (y[36]), .B (n_0_94));
XNOR2_X1 i_0_180 (.ZN (n_0_93), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_179 (.ZN (u[35]), .A (y[35]), .B (n_0_93));
XNOR2_X1 i_0_178 (.ZN (n_0_92), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_177 (.ZN (u[34]), .A (y[34]), .B (n_0_92));
XNOR2_X1 i_0_176 (.ZN (n_0_91), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_175 (.ZN (u[33]), .A (y[33]), .B (n_0_91));
XNOR2_X1 i_0_174 (.ZN (n_0_90), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_173 (.ZN (u[32]), .A (y[32]), .B (n_0_90));
XNOR2_X1 i_0_172 (.ZN (n_0_89), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_171 (.ZN (u[31]), .A (y[31]), .B (n_0_89));
XNOR2_X1 i_0_170 (.ZN (n_0_88), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_169 (.ZN (u[30]), .A (y[30]), .B (n_0_88));
XNOR2_X1 i_0_168 (.ZN (n_0_87), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_167 (.ZN (u[29]), .A (y[29]), .B (n_0_87));
XNOR2_X1 i_0_166 (.ZN (n_0_86), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_165 (.ZN (u[28]), .A (y[28]), .B (n_0_86));
XNOR2_X1 i_0_164 (.ZN (n_0_85), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_163 (.ZN (u[27]), .A (y[27]), .B (n_0_85));
XNOR2_X1 i_0_162 (.ZN (n_0_84), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_161 (.ZN (u[26]), .A (y[26]), .B (n_0_84));
XNOR2_X1 i_0_160 (.ZN (n_0_83), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_159 (.ZN (u[25]), .A (y[25]), .B (n_0_83));
XNOR2_X1 i_0_158 (.ZN (n_0_82), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_157 (.ZN (u[24]), .A (y[24]), .B (n_0_82));
XNOR2_X1 i_0_156 (.ZN (n_0_81), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_155 (.ZN (u[23]), .A (y[23]), .B (n_0_81));
XNOR2_X1 i_0_154 (.ZN (n_0_80), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_153 (.ZN (u[22]), .A (y[22]), .B (n_0_80));
XNOR2_X1 i_0_152 (.ZN (n_0_79), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_151 (.ZN (u[21]), .A (y[21]), .B (n_0_79));
XNOR2_X1 i_0_150 (.ZN (n_0_78), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_149 (.ZN (u[20]), .A (y[20]), .B (n_0_78));
XNOR2_X1 i_0_148 (.ZN (n_0_77), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_147 (.ZN (u[19]), .A (y[19]), .B (n_0_77));
XNOR2_X1 i_0_146 (.ZN (n_0_76), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_145 (.ZN (u[18]), .A (y[18]), .B (n_0_76));
XNOR2_X1 i_0_144 (.ZN (n_0_75), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_143 (.ZN (u[17]), .A (y[17]), .B (n_0_75));
XNOR2_X1 i_0_142 (.ZN (n_0_74), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_141 (.ZN (u[16]), .A (y[16]), .B (n_0_74));
XNOR2_X1 i_0_140 (.ZN (n_0_73), .A (z[15]), .B (x[15]));
XNOR2_X1 i_0_139 (.ZN (u[15]), .A (y[15]), .B (n_0_73));
XNOR2_X1 i_0_138 (.ZN (n_0_72), .A (z[14]), .B (x[14]));
XNOR2_X1 i_0_137 (.ZN (u[14]), .A (y[14]), .B (n_0_72));
XNOR2_X1 i_0_136 (.ZN (n_0_71), .A (z[13]), .B (x[13]));
XNOR2_X2 i_0_135 (.ZN (u[13]), .A (y[13]), .B (n_0_71));
XNOR2_X1 i_0_134 (.ZN (n_0_70), .A (z[12]), .B (x[12]));
XNOR2_X2 i_0_133 (.ZN (u[12]), .A (y[12]), .B (n_0_70));
XNOR2_X2 i_0_132 (.ZN (n_0_69), .A (z[11]), .B (x[11]));
XNOR2_X2 i_0_131 (.ZN (u[11]), .A (y[11]), .B (n_0_69));
NAND2_X2 slo__sro_c12 (.ZN (v[10]), .A1 (n_0_2), .A2 (n_0_3));
XNOR2_X2 i_0_128 (.ZN (n_0_67), .A (x[9]), .B (z[9]));
XNOR2_X2 i_0_127 (.ZN (u[9]), .A (n_0_67), .B (y[9]));
XNOR2_X1 i_0_126 (.ZN (n_0_66), .A (z[8]), .B (x[8]));
XNOR2_X2 i_0_125 (.ZN (u[8]), .A (y[8]), .B (n_0_66));
XOR2_X1 i_0_124 (.Z (u[7]), .A (y[7]), .B (x[7]));
XOR2_X1 i_0_123 (.Z (u[6]), .A (y[6]), .B (x[6]));
NAND2_X2 i_0_122 (.ZN (n_0_65), .A1 (y[63]), .A2 (z[63]));
NOR2_X4 i_0_121 (.ZN (n_0_64), .A1 (y[63]), .A2 (z[63]));
OAI21_X1 i_0_120 (.ZN (v[63]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_121));
OAI21_X1 i_0_119 (.ZN (v[62]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_120));
OAI21_X1 i_0_118 (.ZN (v[61]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_119));
OAI21_X1 i_0_117 (.ZN (v[60]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_118));
OAI21_X1 i_0_116 (.ZN (v[59]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_117));
OAI21_X1 i_0_115 (.ZN (v[58]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_116));
OAI21_X1 i_0_114 (.ZN (v[57]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_115));
OAI21_X1 i_0_113 (.ZN (v[56]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_114));
OAI21_X1 i_0_112 (.ZN (v[55]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_113));
OAI21_X1 i_0_111 (.ZN (v[54]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_112));
OAI21_X1 i_0_110 (.ZN (v[53]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_111));
OAI21_X1 i_0_109 (.ZN (v[52]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_110));
OAI21_X1 i_0_108 (.ZN (v[51]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_109));
OAI21_X1 i_0_107 (.ZN (v[50]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_108));
OAI21_X1 i_0_106 (.ZN (v[49]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_107));
OAI21_X1 i_0_105 (.ZN (v[48]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_106));
OAI21_X1 i_0_104 (.ZN (v[47]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_105));
OAI21_X1 i_0_103 (.ZN (v[46]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_104));
OAI21_X1 i_0_102 (.ZN (v[45]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_103));
OAI21_X1 i_0_101 (.ZN (v[44]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_102));
OAI21_X1 i_0_100 (.ZN (v[43]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_101));
OAI21_X1 i_0_99 (.ZN (v[42]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_100));
OAI21_X1 i_0_98 (.ZN (v[41]), .A (n_0_65), .B1 (n_0_64), .B2 (n_0_99));
NAND2_X1 i_0_97 (.ZN (n_0_63), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_96 (.ZN (n_0_62), .A (y[63]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_95 (.ZN (v[40]), .A1 (n_0_63), .A2 (n_0_62));
NAND2_X1 i_0_94 (.ZN (n_0_61), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_93 (.ZN (n_0_60), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_92 (.ZN (v[39]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_91 (.ZN (n_0_59), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_90 (.ZN (n_0_58), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_89 (.ZN (v[38]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_88 (.ZN (n_0_57), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_87 (.ZN (n_0_56), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_86 (.ZN (v[37]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_85 (.ZN (n_0_55), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_84 (.ZN (n_0_54), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_83 (.ZN (v[36]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_82 (.ZN (n_0_53), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_81 (.ZN (n_0_52), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_80 (.ZN (v[35]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_79 (.ZN (n_0_51), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_78 (.ZN (n_0_50), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_77 (.ZN (v[34]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_76 (.ZN (n_0_49), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_75 (.ZN (n_0_48), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_74 (.ZN (v[33]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_73 (.ZN (n_0_47), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_72 (.ZN (n_0_46), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_71 (.ZN (v[32]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_70 (.ZN (n_0_45), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_69 (.ZN (n_0_44), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_68 (.ZN (v[31]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_67 (.ZN (n_0_43), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_66 (.ZN (n_0_42), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_65 (.ZN (v[30]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_64 (.ZN (n_0_41), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_63 (.ZN (n_0_40), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_62 (.ZN (v[29]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_61 (.ZN (n_0_39), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_60 (.ZN (n_0_38), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_59 (.ZN (v[28]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_58 (.ZN (n_0_37), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_57 (.ZN (n_0_36), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_56 (.ZN (v[27]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_55 (.ZN (n_0_35), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_54 (.ZN (n_0_34), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_53 (.ZN (v[26]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_52 (.ZN (n_0_33), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_51 (.ZN (n_0_32), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_50 (.ZN (v[25]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_49 (.ZN (n_0_31), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_48 (.ZN (n_0_30), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_47 (.ZN (v[24]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_46 (.ZN (n_0_29), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_45 (.ZN (n_0_28), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_44 (.ZN (v[23]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_43 (.ZN (n_0_27), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_42 (.ZN (n_0_26), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_41 (.ZN (v[22]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_40 (.ZN (n_0_25), .A1 (y[20]), .A2 (z[20]));
OAI21_X1 i_0_39 (.ZN (n_0_24), .A (x[20]), .B1 (z[20]), .B2 (y[20]));
NAND2_X1 i_0_38 (.ZN (v[21]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_37 (.ZN (n_0_23), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_36 (.ZN (n_0_22), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_35 (.ZN (v[20]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_34 (.ZN (n_0_21), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_33 (.ZN (n_0_20), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_32 (.ZN (v[19]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_31 (.ZN (n_0_19), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_30 (.ZN (n_0_18), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_29 (.ZN (v[18]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_28 (.ZN (n_0_17), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_27 (.ZN (n_0_16), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_26 (.ZN (v[17]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_25 (.ZN (n_0_15), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_24 (.ZN (n_0_14), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_23 (.ZN (v[16]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_22 (.ZN (n_0_13), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_21 (.ZN (n_0_12), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_20 (.ZN (v[15]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_19 (.ZN (n_0_11), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_18 (.ZN (n_0_10), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X2 i_0_17 (.ZN (v[14]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_16 (.ZN (n_0_9), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_15 (.ZN (n_0_8), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X4 i_0_14 (.ZN (v[13]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_13 (.ZN (n_0_7), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_12 (.ZN (n_0_6), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X4 i_0_11 (.ZN (v[12]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_10 (.ZN (n_0_5), .A1 (z[10]), .A2 (x[10]));
OAI21_X1 i_0_9 (.ZN (n_0_4), .A (y[10]), .B1 (z[10]), .B2 (x[10]));
NAND2_X2 i_0_8 (.ZN (v[11]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_7 (.ZN (n_0_3), .A1 (z[9]), .A2 (x[9]));
OAI21_X1 i_0_6 (.ZN (n_0_2), .A (y[9]), .B1 (z[9]), .B2 (x[9]));
NAND2_X1 i_0_4 (.ZN (n_0_1), .A1 (z[8]), .A2 (x[8]));
OAI21_X1 i_0_3 (.ZN (n_0_0), .A (y[8]), .B1 (z[8]), .B2 (x[8]));
NAND2_X1 i_0_2 (.ZN (v[9]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_1 (.ZN (v[8]), .A1 (y[7]), .A2 (x[7]));
AND2_X1 i_0_0 (.ZN (v[7]), .A1 (y[6]), .A2 (x[6]));
BUF_X2 drc_ipo_c3 (.Z (drc_ipo_n3), .A (n_0_98));
XNOR2_X2 slo__mro_c4 (.ZN (slo__mro_n6), .A (z[10]), .B (x[10]));
XNOR2_X2 slo__mro_c5 (.ZN (u[10]), .A (slo__mro_n6), .B (y[10]));

endmodule //CSA__2_5

module CSA__2_2 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire slo__mro_n7;
wire slo__mro_n8;


XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[63]), .B (x[63]));
XOR2_X1 i_0_158 (.Z (u[63]), .A (z[63]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[38]), .A (z[38]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[37]), .B (x[63]));
XNOR2_X1 i_0_155 (.ZN (u[37]), .A (y[37]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_153 (.ZN (u[36]), .A (y[36]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_151 (.ZN (u[35]), .A (y[35]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_149 (.ZN (u[34]), .A (y[34]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_147 (.ZN (u[33]), .A (y[33]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_145 (.ZN (u[32]), .A (y[32]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_143 (.ZN (u[31]), .A (y[31]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_141 (.ZN (u[30]), .A (y[30]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_139 (.ZN (u[29]), .A (y[29]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_137 (.ZN (u[28]), .A (y[28]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_135 (.ZN (u[27]), .A (y[27]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_133 (.ZN (u[26]), .A (y[26]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_131 (.ZN (u[25]), .A (y[25]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_129 (.ZN (u[24]), .A (y[24]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_127 (.ZN (u[23]), .A (y[23]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_125 (.ZN (u[22]), .A (y[22]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_123 (.ZN (u[21]), .A (y[21]), .B (n_0_76));
XNOR2_X1 i_0_122 (.ZN (n_0_75), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_121 (.ZN (u[20]), .A (y[20]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_119 (.ZN (u[19]), .A (y[19]), .B (n_0_74));
XNOR2_X1 i_0_118 (.ZN (n_0_73), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_117 (.ZN (u[18]), .A (y[18]), .B (n_0_73));
XNOR2_X1 i_0_116 (.ZN (n_0_72), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_115 (.ZN (u[17]), .A (y[17]), .B (n_0_72));
XNOR2_X1 i_0_114 (.ZN (n_0_71), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_113 (.ZN (u[16]), .A (y[16]), .B (n_0_71));
XNOR2_X1 i_0_112 (.ZN (n_0_70), .A (z[15]), .B (x[15]));
XNOR2_X1 i_0_111 (.ZN (u[15]), .A (y[15]), .B (n_0_70));
XNOR2_X1 i_0_110 (.ZN (n_0_69), .A (z[14]), .B (x[14]));
XNOR2_X1 i_0_109 (.ZN (u[14]), .A (y[14]), .B (n_0_69));
XNOR2_X1 i_0_108 (.ZN (n_0_68), .A (z[13]), .B (x[13]));
XNOR2_X2 i_0_107 (.ZN (u[13]), .A (y[13]), .B (n_0_68));
XNOR2_X1 i_0_106 (.ZN (n_0_67), .A (z[12]), .B (x[12]));
XNOR2_X1 i_0_105 (.ZN (u[12]), .A (y[12]), .B (n_0_67));
XNOR2_X2 i_0_104 (.ZN (n_0_66), .A (z[11]), .B (x[11]));
XNOR2_X2 i_0_103 (.ZN (u[11]), .A (y[11]), .B (n_0_66));
XNOR2_X2 i_0_102 (.ZN (n_0_65), .A (z[10]), .B (x[10]));
XNOR2_X2 i_0_101 (.ZN (u[10]), .A (n_0_65), .B (y[10]));
XNOR2_X1 i_0_100 (.ZN (n_0_64), .A (z[9]), .B (x[9]));
XNOR2_X2 i_0_99 (.ZN (u[9]), .A (n_0_64), .B (y[9]));
XNOR2_X1 i_0_98 (.ZN (n_0_63), .A (z[8]), .B (x[8]));
XNOR2_X2 i_0_97 (.ZN (u[8]), .A (y[8]), .B (n_0_63));
XOR2_X1 i_0_96 (.Z (u[7]), .A (y[7]), .B (x[7]));
NAND2_X1 i_0_95 (.ZN (n_0_62), .A1 (y[63]), .A2 (x[63]));
OAI21_X1 i_0_94 (.ZN (n_0_61), .A (z[63]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_93 (.ZN (v[63]), .A1 (n_0_62), .A2 (n_0_61));
OAI21_X1 i_0_92 (.ZN (n_0_60), .A (z[38]), .B1 (x[63]), .B2 (y[63]));
NAND2_X1 i_0_91 (.ZN (v[39]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[37]), .A2 (x[63]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[37]), .B1 (z[37]), .B2 (x[63]));
NAND2_X1 i_0_88 (.ZN (v[38]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_85 (.ZN (v[37]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_82 (.ZN (v[36]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_79 (.ZN (v[35]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_76 (.ZN (v[34]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_73 (.ZN (v[33]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_70 (.ZN (v[32]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_67 (.ZN (v[31]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_64 (.ZN (v[30]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_61 (.ZN (v[29]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_58 (.ZN (v[28]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_55 (.ZN (v[27]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_52 (.ZN (v[26]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_49 (.ZN (v[25]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_46 (.ZN (v[24]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_43 (.ZN (v[23]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_40 (.ZN (v[22]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_37 (.ZN (v[21]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_34 (.ZN (v[20]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_31 (.ZN (v[19]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_28 (.ZN (v[18]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_25 (.ZN (v[17]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_22 (.ZN (v[16]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_19 (.ZN (v[15]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[13]), .A2 (x[13]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[13]), .B1 (z[13]), .B2 (x[13]));
NAND2_X1 i_0_16 (.ZN (v[14]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[12]), .A2 (x[12]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[12]), .B1 (z[12]), .B2 (x[12]));
NAND2_X1 i_0_13 (.ZN (v[13]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[11]), .A2 (x[11]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[11]), .B1 (z[11]), .B2 (x[11]));
NAND2_X1 i_0_10 (.ZN (v[12]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[10]), .A2 (x[10]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[10]), .B1 (z[10]), .B2 (x[10]));
NAND2_X2 i_0_7 (.ZN (v[11]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X2 i_0_6 (.ZN (n_0_3), .A1 (z[9]), .A2 (x[9]));
OAI21_X2 i_0_5 (.ZN (n_0_2), .A (y[9]), .B1 (z[9]), .B2 (x[9]));
NAND2_X4 i_0_4 (.ZN (v[10]), .A1 (n_0_2), .A2 (n_0_3));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[8]), .A2 (x[8]));
AND2_X1 i_0_0 (.ZN (v[8]), .A1 (y[7]), .A2 (x[7]));
OR2_X2 slo__mro_c11 (.ZN (slo__mro_n8), .A1 (x[8]), .A2 (z[8]));
NAND2_X1 slo__mro_c12 (.ZN (slo__mro_n7), .A1 (y[8]), .A2 (slo__mro_n8));
NAND2_X2 slo__mro_c13 (.ZN (v[9]), .A1 (slo__mro_n7), .A2 (n_0_1));

endmodule //CSA__2_2

module CSA__0_69 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;


XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[62]), .B (x[62]));
XOR2_X1 i_0_158 (.Z (u[63]), .A (z[62]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[44]), .A (z[44]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[43]), .B (x[62]));
XNOR2_X1 i_0_155 (.ZN (u[43]), .A (y[43]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_153 (.ZN (u[42]), .A (y[42]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_151 (.ZN (u[41]), .A (y[41]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_149 (.ZN (u[40]), .A (y[40]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_147 (.ZN (u[39]), .A (y[39]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_145 (.ZN (u[38]), .A (y[38]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_143 (.ZN (u[37]), .A (y[37]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_141 (.ZN (u[36]), .A (y[36]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_139 (.ZN (u[35]), .A (y[35]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_137 (.ZN (u[34]), .A (y[34]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_135 (.ZN (u[33]), .A (y[33]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_133 (.ZN (u[32]), .A (y[32]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_131 (.ZN (u[31]), .A (y[31]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_129 (.ZN (u[30]), .A (y[30]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_127 (.ZN (u[29]), .A (y[29]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_125 (.ZN (u[28]), .A (y[28]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_123 (.ZN (u[27]), .A (y[27]), .B (n_0_76));
XNOR2_X1 i_0_122 (.ZN (n_0_75), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_121 (.ZN (u[26]), .A (y[26]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_119 (.ZN (u[25]), .A (y[25]), .B (n_0_74));
XNOR2_X1 i_0_118 (.ZN (n_0_73), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_117 (.ZN (u[24]), .A (y[24]), .B (n_0_73));
XNOR2_X1 i_0_116 (.ZN (n_0_72), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_115 (.ZN (u[23]), .A (y[23]), .B (n_0_72));
XNOR2_X1 i_0_114 (.ZN (n_0_71), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_113 (.ZN (u[22]), .A (y[22]), .B (n_0_71));
XNOR2_X1 i_0_112 (.ZN (n_0_70), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_111 (.ZN (u[21]), .A (y[21]), .B (n_0_70));
XNOR2_X1 i_0_110 (.ZN (n_0_69), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_109 (.ZN (u[20]), .A (y[20]), .B (n_0_69));
XNOR2_X1 i_0_108 (.ZN (n_0_68), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_107 (.ZN (u[19]), .A (y[19]), .B (n_0_68));
XNOR2_X1 i_0_106 (.ZN (n_0_67), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_105 (.ZN (u[18]), .A (y[18]), .B (n_0_67));
XNOR2_X1 i_0_104 (.ZN (n_0_66), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_103 (.ZN (u[17]), .A (y[17]), .B (n_0_66));
XNOR2_X2 i_0_102 (.ZN (n_0_65), .A (z[16]), .B (x[16]));
XNOR2_X1 i_0_101 (.ZN (u[16]), .A (y[16]), .B (n_0_65));
XNOR2_X1 i_0_100 (.ZN (n_0_64), .A (z[15]), .B (x[15]));
XNOR2_X2 i_0_99 (.ZN (u[15]), .A (y[15]), .B (n_0_64));
XNOR2_X1 i_0_98 (.ZN (n_0_63), .A (z[14]), .B (x[14]));
XNOR2_X2 i_0_97 (.ZN (u[14]), .A (y[14]), .B (n_0_63));
XOR2_X2 i_0_96 (.Z (u[13]), .A (y[13]), .B (x[13]));
NOR2_X1 i_0_95 (.ZN (n_0_62), .A1 (y[62]), .A2 (x[62]));
AOI21_X1 i_0_94 (.ZN (n_0_61), .A (z[62]), .B1 (x[62]), .B2 (y[62]));
NOR2_X1 i_0_93 (.ZN (v[63]), .A1 (n_0_62), .A2 (n_0_61));
AOI21_X1 i_0_92 (.ZN (n_0_60), .A (z[44]), .B1 (x[62]), .B2 (y[62]));
NOR2_X1 i_0_91 (.ZN (v[45]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[43]), .A2 (x[62]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[43]), .B1 (z[43]), .B2 (x[62]));
NAND2_X1 i_0_88 (.ZN (v[44]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_85 (.ZN (v[43]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_82 (.ZN (v[42]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_79 (.ZN (v[41]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_76 (.ZN (v[40]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_73 (.ZN (v[39]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_70 (.ZN (v[38]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_67 (.ZN (v[37]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_64 (.ZN (v[36]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_61 (.ZN (v[35]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_58 (.ZN (v[34]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_55 (.ZN (v[33]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_52 (.ZN (v[32]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_49 (.ZN (v[31]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_46 (.ZN (v[30]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_43 (.ZN (v[29]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_40 (.ZN (v[28]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_37 (.ZN (v[27]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_34 (.ZN (v[26]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_31 (.ZN (v[25]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_28 (.ZN (v[24]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_25 (.ZN (v[23]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_22 (.ZN (v[22]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_19 (.ZN (v[21]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_16 (.ZN (v[20]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_13 (.ZN (v[19]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_10 (.ZN (v[18]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[16]), .A2 (x[16]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[16]), .B1 (z[16]), .B2 (x[16]));
NAND2_X1 i_0_7 (.ZN (v[17]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[15]), .A2 (x[15]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[15]), .B1 (z[15]), .B2 (x[15]));
NAND2_X1 i_0_4 (.ZN (v[16]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[14]), .A2 (x[14]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[14]), .B1 (z[14]), .B2 (x[14]));
NAND2_X1 i_0_1 (.ZN (v[15]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[14]), .A1 (y[13]), .A2 (x[13]));

endmodule //CSA__0_69

module CSA__1_5 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;


XOR2_X1 i_0_159 (.Z (n_0_93), .A (y[62]), .B (x[62]));
XOR2_X1 i_0_158 (.Z (u[63]), .A (z[62]), .B (n_0_93));
XOR2_X1 i_0_157 (.Z (u[47]), .A (z[47]), .B (n_0_93));
XNOR2_X1 i_0_156 (.ZN (n_0_92), .A (z[46]), .B (x[62]));
XNOR2_X1 i_0_155 (.ZN (u[46]), .A (y[46]), .B (n_0_92));
XNOR2_X1 i_0_154 (.ZN (n_0_91), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_153 (.ZN (u[45]), .A (y[45]), .B (n_0_91));
XNOR2_X1 i_0_152 (.ZN (n_0_90), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_151 (.ZN (u[44]), .A (y[44]), .B (n_0_90));
XNOR2_X1 i_0_150 (.ZN (n_0_89), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_149 (.ZN (u[43]), .A (y[43]), .B (n_0_89));
XNOR2_X1 i_0_148 (.ZN (n_0_88), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_147 (.ZN (u[42]), .A (y[42]), .B (n_0_88));
XNOR2_X1 i_0_146 (.ZN (n_0_87), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_145 (.ZN (u[41]), .A (y[41]), .B (n_0_87));
XNOR2_X1 i_0_144 (.ZN (n_0_86), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_143 (.ZN (u[40]), .A (y[40]), .B (n_0_86));
XNOR2_X1 i_0_142 (.ZN (n_0_85), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_141 (.ZN (u[39]), .A (y[39]), .B (n_0_85));
XNOR2_X1 i_0_140 (.ZN (n_0_84), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_139 (.ZN (u[38]), .A (y[38]), .B (n_0_84));
XNOR2_X1 i_0_138 (.ZN (n_0_83), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_137 (.ZN (u[37]), .A (y[37]), .B (n_0_83));
XNOR2_X1 i_0_136 (.ZN (n_0_82), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_135 (.ZN (u[36]), .A (y[36]), .B (n_0_82));
XNOR2_X1 i_0_134 (.ZN (n_0_81), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_133 (.ZN (u[35]), .A (y[35]), .B (n_0_81));
XNOR2_X1 i_0_132 (.ZN (n_0_80), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_131 (.ZN (u[34]), .A (y[34]), .B (n_0_80));
XNOR2_X1 i_0_130 (.ZN (n_0_79), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_129 (.ZN (u[33]), .A (y[33]), .B (n_0_79));
XNOR2_X1 i_0_128 (.ZN (n_0_78), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_127 (.ZN (u[32]), .A (y[32]), .B (n_0_78));
XNOR2_X1 i_0_126 (.ZN (n_0_77), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_125 (.ZN (u[31]), .A (y[31]), .B (n_0_77));
XNOR2_X1 i_0_124 (.ZN (n_0_76), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_123 (.ZN (u[30]), .A (y[30]), .B (n_0_76));
XNOR2_X1 i_0_122 (.ZN (n_0_75), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_121 (.ZN (u[29]), .A (y[29]), .B (n_0_75));
XNOR2_X1 i_0_120 (.ZN (n_0_74), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_119 (.ZN (u[28]), .A (y[28]), .B (n_0_74));
XNOR2_X1 i_0_118 (.ZN (n_0_73), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_117 (.ZN (u[27]), .A (y[27]), .B (n_0_73));
XNOR2_X1 i_0_116 (.ZN (n_0_72), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_115 (.ZN (u[26]), .A (y[26]), .B (n_0_72));
XNOR2_X1 i_0_114 (.ZN (n_0_71), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_113 (.ZN (u[25]), .A (y[25]), .B (n_0_71));
XNOR2_X1 i_0_112 (.ZN (n_0_70), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_111 (.ZN (u[24]), .A (y[24]), .B (n_0_70));
XNOR2_X1 i_0_110 (.ZN (n_0_69), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_109 (.ZN (u[23]), .A (y[23]), .B (n_0_69));
XNOR2_X1 i_0_108 (.ZN (n_0_68), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_107 (.ZN (u[22]), .A (y[22]), .B (n_0_68));
XNOR2_X1 i_0_106 (.ZN (n_0_67), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_105 (.ZN (u[21]), .A (y[21]), .B (n_0_67));
XNOR2_X1 i_0_104 (.ZN (n_0_66), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_103 (.ZN (u[20]), .A (y[20]), .B (n_0_66));
XNOR2_X1 i_0_102 (.ZN (n_0_65), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_101 (.ZN (u[19]), .A (y[19]), .B (n_0_65));
XNOR2_X1 i_0_100 (.ZN (n_0_64), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_99 (.ZN (u[18]), .A (y[18]), .B (n_0_64));
XNOR2_X1 i_0_98 (.ZN (n_0_63), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_97 (.ZN (u[17]), .A (y[17]), .B (n_0_63));
XOR2_X1 i_0_96 (.Z (u[16]), .A (y[16]), .B (x[16]));
NOR2_X1 i_0_95 (.ZN (n_0_62), .A1 (y[62]), .A2 (x[62]));
AOI21_X1 i_0_94 (.ZN (n_0_61), .A (z[62]), .B1 (x[62]), .B2 (y[62]));
NOR2_X1 i_0_93 (.ZN (v[63]), .A1 (n_0_62), .A2 (n_0_61));
AOI21_X1 i_0_92 (.ZN (n_0_60), .A (z[47]), .B1 (x[62]), .B2 (y[62]));
NOR2_X1 i_0_91 (.ZN (v[48]), .A1 (n_0_62), .A2 (n_0_60));
NAND2_X1 i_0_90 (.ZN (n_0_59), .A1 (z[46]), .A2 (x[62]));
OAI21_X1 i_0_89 (.ZN (n_0_58), .A (y[46]), .B1 (z[46]), .B2 (x[62]));
NAND2_X1 i_0_88 (.ZN (v[47]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_87 (.ZN (n_0_57), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_86 (.ZN (n_0_56), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_85 (.ZN (v[46]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_84 (.ZN (n_0_55), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_83 (.ZN (n_0_54), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_82 (.ZN (v[45]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_81 (.ZN (n_0_53), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_80 (.ZN (n_0_52), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_79 (.ZN (v[44]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_78 (.ZN (n_0_51), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_77 (.ZN (n_0_50), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_76 (.ZN (v[43]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_75 (.ZN (n_0_49), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_74 (.ZN (n_0_48), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_73 (.ZN (v[42]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_72 (.ZN (n_0_47), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_71 (.ZN (n_0_46), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_70 (.ZN (v[41]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_69 (.ZN (n_0_45), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_68 (.ZN (n_0_44), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_67 (.ZN (v[40]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_66 (.ZN (n_0_43), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_65 (.ZN (n_0_42), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_64 (.ZN (v[39]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_63 (.ZN (n_0_41), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_62 (.ZN (n_0_40), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_61 (.ZN (v[38]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_60 (.ZN (n_0_39), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_59 (.ZN (n_0_38), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_58 (.ZN (v[37]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_57 (.ZN (n_0_37), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_56 (.ZN (n_0_36), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_55 (.ZN (v[36]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_54 (.ZN (n_0_35), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_53 (.ZN (n_0_34), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_52 (.ZN (v[35]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_51 (.ZN (n_0_33), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_50 (.ZN (n_0_32), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_49 (.ZN (v[34]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_48 (.ZN (n_0_31), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_47 (.ZN (n_0_30), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_46 (.ZN (v[33]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_45 (.ZN (n_0_29), .A1 (z[31]), .A2 (x[31]));
OAI21_X1 i_0_44 (.ZN (n_0_28), .A (y[31]), .B1 (z[31]), .B2 (x[31]));
NAND2_X1 i_0_43 (.ZN (v[32]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_42 (.ZN (n_0_27), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_41 (.ZN (n_0_26), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_40 (.ZN (v[31]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_39 (.ZN (n_0_25), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_38 (.ZN (n_0_24), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_37 (.ZN (v[30]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_36 (.ZN (n_0_23), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_35 (.ZN (n_0_22), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_34 (.ZN (v[29]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_33 (.ZN (n_0_21), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_32 (.ZN (n_0_20), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_31 (.ZN (v[28]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_30 (.ZN (n_0_19), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_29 (.ZN (n_0_18), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_28 (.ZN (v[27]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_27 (.ZN (n_0_17), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_26 (.ZN (n_0_16), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_25 (.ZN (v[26]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_24 (.ZN (n_0_15), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_23 (.ZN (n_0_14), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_22 (.ZN (v[25]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_21 (.ZN (n_0_13), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_20 (.ZN (n_0_12), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_19 (.ZN (v[24]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_18 (.ZN (n_0_11), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_17 (.ZN (n_0_10), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_16 (.ZN (v[23]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_15 (.ZN (n_0_9), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_14 (.ZN (n_0_8), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_13 (.ZN (v[22]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_11 (.ZN (n_0_6), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_10 (.ZN (v[21]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_9 (.ZN (n_0_5), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_8 (.ZN (n_0_4), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_7 (.ZN (v[20]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_6 (.ZN (n_0_3), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_5 (.ZN (n_0_2), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_4 (.ZN (v[19]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_3 (.ZN (n_0_1), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_2 (.ZN (n_0_0), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_1 (.ZN (v[18]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_0 (.ZN (v[17]), .A1 (y[16]), .A2 (x[16]));

endmodule //CSA__1_5

module CSA__1_2 (x, y, z, u, v);

output [63:0] u;
output [63:0] v;
input [63:0] x;
input [63:0] y;
input [63:0] z;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;


XOR2_X1 i_0_166 (.Z (n_0_96), .A (y[63]), .B (x[63]));
XOR2_X1 i_0_165 (.Z (u[63]), .A (z[63]), .B (n_0_96));
XOR2_X1 i_0_164 (.Z (u[48]), .A (z[48]), .B (n_0_96));
XNOR2_X1 i_0_163 (.ZN (n_0_95), .A (z[47]), .B (x[63]));
XNOR2_X1 i_0_162 (.ZN (u[47]), .A (y[47]), .B (n_0_95));
XNOR2_X1 i_0_161 (.ZN (n_0_94), .A (z[46]), .B (x[63]));
XNOR2_X1 i_0_160 (.ZN (u[46]), .A (y[46]), .B (n_0_94));
XNOR2_X1 i_0_159 (.ZN (n_0_93), .A (z[45]), .B (x[45]));
XNOR2_X1 i_0_158 (.ZN (u[45]), .A (y[45]), .B (n_0_93));
XNOR2_X1 i_0_157 (.ZN (n_0_92), .A (z[44]), .B (x[44]));
XNOR2_X1 i_0_156 (.ZN (u[44]), .A (y[44]), .B (n_0_92));
XNOR2_X1 i_0_155 (.ZN (n_0_91), .A (z[43]), .B (x[43]));
XNOR2_X1 i_0_154 (.ZN (u[43]), .A (y[43]), .B (n_0_91));
XNOR2_X1 i_0_153 (.ZN (n_0_90), .A (z[42]), .B (x[42]));
XNOR2_X1 i_0_152 (.ZN (u[42]), .A (y[42]), .B (n_0_90));
XNOR2_X1 i_0_151 (.ZN (n_0_89), .A (z[41]), .B (x[41]));
XNOR2_X1 i_0_150 (.ZN (u[41]), .A (y[41]), .B (n_0_89));
XNOR2_X1 i_0_149 (.ZN (n_0_88), .A (z[40]), .B (x[40]));
XNOR2_X1 i_0_148 (.ZN (u[40]), .A (y[40]), .B (n_0_88));
XNOR2_X1 i_0_147 (.ZN (n_0_87), .A (z[39]), .B (x[39]));
XNOR2_X1 i_0_146 (.ZN (u[39]), .A (y[39]), .B (n_0_87));
XNOR2_X1 i_0_145 (.ZN (n_0_86), .A (z[38]), .B (x[38]));
XNOR2_X1 i_0_144 (.ZN (u[38]), .A (y[38]), .B (n_0_86));
XNOR2_X1 i_0_143 (.ZN (n_0_85), .A (z[37]), .B (x[37]));
XNOR2_X1 i_0_142 (.ZN (u[37]), .A (y[37]), .B (n_0_85));
XNOR2_X1 i_0_141 (.ZN (n_0_84), .A (z[36]), .B (x[36]));
XNOR2_X1 i_0_140 (.ZN (u[36]), .A (y[36]), .B (n_0_84));
XNOR2_X1 i_0_139 (.ZN (n_0_83), .A (z[35]), .B (x[35]));
XNOR2_X1 i_0_138 (.ZN (u[35]), .A (y[35]), .B (n_0_83));
XNOR2_X1 i_0_137 (.ZN (n_0_82), .A (z[34]), .B (x[34]));
XNOR2_X1 i_0_136 (.ZN (u[34]), .A (y[34]), .B (n_0_82));
XNOR2_X1 i_0_135 (.ZN (n_0_81), .A (z[33]), .B (x[33]));
XNOR2_X1 i_0_134 (.ZN (u[33]), .A (y[33]), .B (n_0_81));
XNOR2_X1 i_0_133 (.ZN (n_0_80), .A (z[32]), .B (x[32]));
XNOR2_X1 i_0_132 (.ZN (u[32]), .A (y[32]), .B (n_0_80));
XNOR2_X1 i_0_131 (.ZN (n_0_79), .A (z[31]), .B (x[31]));
XNOR2_X1 i_0_130 (.ZN (u[31]), .A (y[31]), .B (n_0_79));
XNOR2_X1 i_0_129 (.ZN (n_0_78), .A (z[30]), .B (x[30]));
XNOR2_X1 i_0_128 (.ZN (u[30]), .A (y[30]), .B (n_0_78));
XNOR2_X1 i_0_127 (.ZN (n_0_77), .A (z[29]), .B (x[29]));
XNOR2_X1 i_0_126 (.ZN (u[29]), .A (y[29]), .B (n_0_77));
XNOR2_X1 i_0_125 (.ZN (n_0_76), .A (z[28]), .B (x[28]));
XNOR2_X1 i_0_124 (.ZN (u[28]), .A (y[28]), .B (n_0_76));
XNOR2_X1 i_0_123 (.ZN (n_0_75), .A (z[27]), .B (x[27]));
XNOR2_X1 i_0_122 (.ZN (u[27]), .A (y[27]), .B (n_0_75));
XNOR2_X1 i_0_121 (.ZN (n_0_74), .A (z[26]), .B (x[26]));
XNOR2_X1 i_0_120 (.ZN (u[26]), .A (y[26]), .B (n_0_74));
XNOR2_X1 i_0_119 (.ZN (n_0_73), .A (z[25]), .B (x[25]));
XNOR2_X1 i_0_118 (.ZN (u[25]), .A (y[25]), .B (n_0_73));
XNOR2_X1 i_0_117 (.ZN (n_0_72), .A (z[24]), .B (x[24]));
XNOR2_X1 i_0_116 (.ZN (u[24]), .A (y[24]), .B (n_0_72));
XNOR2_X1 i_0_115 (.ZN (n_0_71), .A (z[23]), .B (x[23]));
XNOR2_X1 i_0_114 (.ZN (u[23]), .A (y[23]), .B (n_0_71));
XNOR2_X1 i_0_113 (.ZN (n_0_70), .A (z[22]), .B (x[22]));
XNOR2_X1 i_0_112 (.ZN (u[22]), .A (y[22]), .B (n_0_70));
XNOR2_X1 i_0_111 (.ZN (n_0_69), .A (z[21]), .B (x[21]));
XNOR2_X1 i_0_110 (.ZN (u[21]), .A (y[21]), .B (n_0_69));
XNOR2_X1 i_0_109 (.ZN (n_0_68), .A (z[20]), .B (x[20]));
XNOR2_X1 i_0_108 (.ZN (u[20]), .A (y[20]), .B (n_0_68));
XNOR2_X1 i_0_107 (.ZN (n_0_67), .A (z[19]), .B (x[19]));
XNOR2_X1 i_0_106 (.ZN (u[19]), .A (y[19]), .B (n_0_67));
XNOR2_X1 i_0_105 (.ZN (n_0_66), .A (z[18]), .B (x[18]));
XNOR2_X1 i_0_104 (.ZN (u[18]), .A (y[18]), .B (n_0_66));
XNOR2_X1 i_0_103 (.ZN (n_0_65), .A (z[17]), .B (x[17]));
XNOR2_X1 i_0_102 (.ZN (u[17]), .A (y[17]), .B (n_0_65));
XOR2_X1 i_0_101 (.Z (u[16]), .A (y[16]), .B (x[16]));
XOR2_X1 i_0_100 (.Z (u[15]), .A (y[15]), .B (x[15]));
NOR2_X1 i_0_99 (.ZN (n_0_64), .A1 (y[63]), .A2 (x[63]));
AOI21_X1 i_0_98 (.ZN (n_0_63), .A (z[63]), .B1 (x[63]), .B2 (y[63]));
NOR2_X1 i_0_97 (.ZN (v[63]), .A1 (n_0_64), .A2 (n_0_63));
AOI21_X1 i_0_96 (.ZN (n_0_62), .A (z[48]), .B1 (x[63]), .B2 (y[63]));
NOR2_X1 i_0_95 (.ZN (v[49]), .A1 (n_0_64), .A2 (n_0_62));
NAND2_X1 i_0_94 (.ZN (n_0_61), .A1 (z[47]), .A2 (x[63]));
OAI21_X1 i_0_93 (.ZN (n_0_60), .A (y[47]), .B1 (z[47]), .B2 (x[63]));
NAND2_X1 i_0_92 (.ZN (v[48]), .A1 (n_0_61), .A2 (n_0_60));
NAND2_X1 i_0_91 (.ZN (n_0_59), .A1 (z[46]), .A2 (x[63]));
OAI21_X1 i_0_90 (.ZN (n_0_58), .A (y[46]), .B1 (z[46]), .B2 (x[63]));
NAND2_X1 i_0_89 (.ZN (v[47]), .A1 (n_0_59), .A2 (n_0_58));
NAND2_X1 i_0_88 (.ZN (n_0_57), .A1 (z[45]), .A2 (x[45]));
OAI21_X1 i_0_87 (.ZN (n_0_56), .A (y[45]), .B1 (z[45]), .B2 (x[45]));
NAND2_X1 i_0_86 (.ZN (v[46]), .A1 (n_0_57), .A2 (n_0_56));
NAND2_X1 i_0_85 (.ZN (n_0_55), .A1 (z[44]), .A2 (x[44]));
OAI21_X1 i_0_84 (.ZN (n_0_54), .A (y[44]), .B1 (z[44]), .B2 (x[44]));
NAND2_X1 i_0_83 (.ZN (v[45]), .A1 (n_0_55), .A2 (n_0_54));
NAND2_X1 i_0_82 (.ZN (n_0_53), .A1 (z[43]), .A2 (x[43]));
OAI21_X1 i_0_81 (.ZN (n_0_52), .A (y[43]), .B1 (z[43]), .B2 (x[43]));
NAND2_X1 i_0_80 (.ZN (v[44]), .A1 (n_0_53), .A2 (n_0_52));
NAND2_X1 i_0_79 (.ZN (n_0_51), .A1 (z[42]), .A2 (x[42]));
OAI21_X1 i_0_78 (.ZN (n_0_50), .A (y[42]), .B1 (z[42]), .B2 (x[42]));
NAND2_X1 i_0_77 (.ZN (v[43]), .A1 (n_0_51), .A2 (n_0_50));
NAND2_X1 i_0_76 (.ZN (n_0_49), .A1 (z[41]), .A2 (x[41]));
OAI21_X1 i_0_75 (.ZN (n_0_48), .A (y[41]), .B1 (z[41]), .B2 (x[41]));
NAND2_X1 i_0_74 (.ZN (v[42]), .A1 (n_0_49), .A2 (n_0_48));
NAND2_X1 i_0_73 (.ZN (n_0_47), .A1 (z[40]), .A2 (x[40]));
OAI21_X1 i_0_72 (.ZN (n_0_46), .A (y[40]), .B1 (z[40]), .B2 (x[40]));
NAND2_X1 i_0_71 (.ZN (v[41]), .A1 (n_0_47), .A2 (n_0_46));
NAND2_X1 i_0_70 (.ZN (n_0_45), .A1 (z[39]), .A2 (x[39]));
OAI21_X1 i_0_69 (.ZN (n_0_44), .A (y[39]), .B1 (z[39]), .B2 (x[39]));
NAND2_X1 i_0_68 (.ZN (v[40]), .A1 (n_0_45), .A2 (n_0_44));
NAND2_X1 i_0_67 (.ZN (n_0_43), .A1 (z[38]), .A2 (x[38]));
OAI21_X1 i_0_66 (.ZN (n_0_42), .A (y[38]), .B1 (z[38]), .B2 (x[38]));
NAND2_X1 i_0_65 (.ZN (v[39]), .A1 (n_0_43), .A2 (n_0_42));
NAND2_X1 i_0_64 (.ZN (n_0_41), .A1 (z[37]), .A2 (x[37]));
OAI21_X1 i_0_63 (.ZN (n_0_40), .A (y[37]), .B1 (z[37]), .B2 (x[37]));
NAND2_X1 i_0_62 (.ZN (v[38]), .A1 (n_0_41), .A2 (n_0_40));
NAND2_X1 i_0_61 (.ZN (n_0_39), .A1 (z[36]), .A2 (x[36]));
OAI21_X1 i_0_60 (.ZN (n_0_38), .A (y[36]), .B1 (z[36]), .B2 (x[36]));
NAND2_X1 i_0_59 (.ZN (v[37]), .A1 (n_0_39), .A2 (n_0_38));
NAND2_X1 i_0_58 (.ZN (n_0_37), .A1 (z[35]), .A2 (x[35]));
OAI21_X1 i_0_57 (.ZN (n_0_36), .A (y[35]), .B1 (z[35]), .B2 (x[35]));
NAND2_X1 i_0_56 (.ZN (v[36]), .A1 (n_0_37), .A2 (n_0_36));
NAND2_X1 i_0_55 (.ZN (n_0_35), .A1 (z[34]), .A2 (x[34]));
OAI21_X1 i_0_54 (.ZN (n_0_34), .A (y[34]), .B1 (z[34]), .B2 (x[34]));
NAND2_X1 i_0_53 (.ZN (v[35]), .A1 (n_0_35), .A2 (n_0_34));
NAND2_X1 i_0_52 (.ZN (n_0_33), .A1 (z[33]), .A2 (x[33]));
OAI21_X1 i_0_51 (.ZN (n_0_32), .A (y[33]), .B1 (z[33]), .B2 (x[33]));
NAND2_X1 i_0_50 (.ZN (v[34]), .A1 (n_0_33), .A2 (n_0_32));
NAND2_X1 i_0_49 (.ZN (n_0_31), .A1 (z[32]), .A2 (x[32]));
OAI21_X1 i_0_48 (.ZN (n_0_30), .A (y[32]), .B1 (z[32]), .B2 (x[32]));
NAND2_X1 i_0_47 (.ZN (v[33]), .A1 (n_0_31), .A2 (n_0_30));
NAND2_X1 i_0_46 (.ZN (n_0_29), .A1 (y[31]), .A2 (z[31]));
OAI21_X1 i_0_45 (.ZN (n_0_28), .A (x[31]), .B1 (z[31]), .B2 (y[31]));
NAND2_X1 i_0_44 (.ZN (v[32]), .A1 (n_0_29), .A2 (n_0_28));
NAND2_X1 i_0_43 (.ZN (n_0_27), .A1 (z[30]), .A2 (x[30]));
OAI21_X1 i_0_42 (.ZN (n_0_26), .A (y[30]), .B1 (z[30]), .B2 (x[30]));
NAND2_X1 i_0_41 (.ZN (v[31]), .A1 (n_0_27), .A2 (n_0_26));
NAND2_X1 i_0_40 (.ZN (n_0_25), .A1 (z[29]), .A2 (x[29]));
OAI21_X1 i_0_39 (.ZN (n_0_24), .A (y[29]), .B1 (z[29]), .B2 (x[29]));
NAND2_X1 i_0_38 (.ZN (v[30]), .A1 (n_0_25), .A2 (n_0_24));
NAND2_X1 i_0_37 (.ZN (n_0_23), .A1 (z[28]), .A2 (x[28]));
OAI21_X1 i_0_36 (.ZN (n_0_22), .A (y[28]), .B1 (z[28]), .B2 (x[28]));
NAND2_X1 i_0_35 (.ZN (v[29]), .A1 (n_0_23), .A2 (n_0_22));
NAND2_X1 i_0_34 (.ZN (n_0_21), .A1 (z[27]), .A2 (x[27]));
OAI21_X1 i_0_33 (.ZN (n_0_20), .A (y[27]), .B1 (z[27]), .B2 (x[27]));
NAND2_X1 i_0_32 (.ZN (v[28]), .A1 (n_0_21), .A2 (n_0_20));
NAND2_X1 i_0_31 (.ZN (n_0_19), .A1 (z[26]), .A2 (x[26]));
OAI21_X1 i_0_30 (.ZN (n_0_18), .A (y[26]), .B1 (z[26]), .B2 (x[26]));
NAND2_X1 i_0_29 (.ZN (v[27]), .A1 (n_0_19), .A2 (n_0_18));
NAND2_X1 i_0_28 (.ZN (n_0_17), .A1 (z[25]), .A2 (x[25]));
OAI21_X1 i_0_27 (.ZN (n_0_16), .A (y[25]), .B1 (z[25]), .B2 (x[25]));
NAND2_X1 i_0_26 (.ZN (v[26]), .A1 (n_0_17), .A2 (n_0_16));
NAND2_X1 i_0_25 (.ZN (n_0_15), .A1 (z[24]), .A2 (x[24]));
OAI21_X1 i_0_24 (.ZN (n_0_14), .A (y[24]), .B1 (z[24]), .B2 (x[24]));
NAND2_X1 i_0_23 (.ZN (v[25]), .A1 (n_0_15), .A2 (n_0_14));
NAND2_X1 i_0_22 (.ZN (n_0_13), .A1 (z[23]), .A2 (x[23]));
OAI21_X1 i_0_21 (.ZN (n_0_12), .A (y[23]), .B1 (z[23]), .B2 (x[23]));
NAND2_X1 i_0_20 (.ZN (v[24]), .A1 (n_0_13), .A2 (n_0_12));
NAND2_X1 i_0_19 (.ZN (n_0_11), .A1 (z[22]), .A2 (x[22]));
OAI21_X1 i_0_18 (.ZN (n_0_10), .A (y[22]), .B1 (z[22]), .B2 (x[22]));
NAND2_X1 i_0_17 (.ZN (v[23]), .A1 (n_0_11), .A2 (n_0_10));
NAND2_X1 i_0_16 (.ZN (n_0_9), .A1 (z[21]), .A2 (x[21]));
OAI21_X1 i_0_15 (.ZN (n_0_8), .A (y[21]), .B1 (z[21]), .B2 (x[21]));
NAND2_X1 i_0_14 (.ZN (v[22]), .A1 (n_0_9), .A2 (n_0_8));
NAND2_X1 i_0_13 (.ZN (n_0_7), .A1 (z[20]), .A2 (x[20]));
OAI21_X1 i_0_12 (.ZN (n_0_6), .A (y[20]), .B1 (z[20]), .B2 (x[20]));
NAND2_X1 i_0_11 (.ZN (v[21]), .A1 (n_0_7), .A2 (n_0_6));
NAND2_X1 i_0_10 (.ZN (n_0_5), .A1 (z[19]), .A2 (x[19]));
OAI21_X1 i_0_9 (.ZN (n_0_4), .A (y[19]), .B1 (z[19]), .B2 (x[19]));
NAND2_X1 i_0_8 (.ZN (v[20]), .A1 (n_0_5), .A2 (n_0_4));
NAND2_X1 i_0_7 (.ZN (n_0_3), .A1 (z[18]), .A2 (x[18]));
OAI21_X1 i_0_6 (.ZN (n_0_2), .A (y[18]), .B1 (z[18]), .B2 (x[18]));
NAND2_X1 i_0_5 (.ZN (v[19]), .A1 (n_0_3), .A2 (n_0_2));
NAND2_X1 i_0_4 (.ZN (n_0_1), .A1 (z[17]), .A2 (x[17]));
OAI21_X1 i_0_3 (.ZN (n_0_0), .A (y[17]), .B1 (z[17]), .B2 (x[17]));
NAND2_X1 i_0_2 (.ZN (v[18]), .A1 (n_0_1), .A2 (n_0_0));
AND2_X1 i_0_1 (.ZN (v[17]), .A1 (y[16]), .A2 (x[16]));
AND2_X1 i_0_0 (.ZN (v[16]), .A1 (y[15]), .A2 (x[15]));

endmodule //CSA__1_2

module products (x, y, \pp[32] , \pp[31] , \pp[30] , \pp[29] , \pp[28] , \pp[27] , 
    \pp[26] , \pp[25] , \pp[24] , \pp[23] , \pp[22] , \pp[21] , \pp[20] , \pp[19] , 
    \pp[18] , \pp[17] , \pp[16] , \pp[15] , \pp[14] , \pp[13] , \pp[12] , \pp[11] , 
    \pp[10] , \pp[9] , \pp[8] , \pp[7] , \pp[6] , \pp[5] , \pp[4] , \pp[3] , \pp[2] , 
    \pp[1] , \pp[0] );

output [63:0] \pp[0] ;
output [63:0] \pp[10] ;
output [63:0] \pp[11] ;
output [63:0] \pp[12] ;
output [63:0] \pp[13] ;
output [63:0] \pp[14] ;
output [63:0] \pp[15] ;
output [63:0] \pp[16] ;
output [63:0] \pp[17] ;
output [63:0] \pp[18] ;
output [63:0] \pp[19] ;
output [63:0] \pp[1] ;
output [63:0] \pp[20] ;
output [63:0] \pp[21] ;
output [63:0] \pp[22] ;
output [63:0] \pp[23] ;
output [63:0] \pp[24] ;
output [63:0] \pp[25] ;
output [63:0] \pp[26] ;
output [63:0] \pp[27] ;
output [63:0] \pp[28] ;
output [63:0] \pp[29] ;
output [63:0] \pp[2] ;
output [63:0] \pp[30] ;
output [63:0] \pp[31] ;
output [63:0] \pp[32] ;
output [63:0] \pp[3] ;
output [63:0] \pp[4] ;
output [63:0] \pp[5] ;
output [63:0] \pp[6] ;
output [63:0] \pp[7] ;
output [63:0] \pp[8] ;
output [63:0] \pp[9] ;
input [31:0] x;
input [31:0] y;
wire slo___n552;
wire slo___n701;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_56;
wire n_0_63;
wire n_0_62;
wire n_0_61;
wire n_0_60;
wire n_0_59;
wire n_0_58;
wire n_0_57;
wire n_0_55;
wire n_0_13;
wire n_0_12;
wire n_0_11;
wire n_0_10;
wire n_0_9;
wire n_0_8;
wire n_0_7;
wire n_0_6;
wire n_0_5;
wire n_0_4;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire sgo__n150;
wire sgo__n157;
wire sgo__n162;
wire sgo__n167;
wire sgo__n172;
wire sgo__n177;
wire sgo__n184;
wire sgo__n205;
wire sgo__n240;
wire sgo__n272;
wire sgo__n301;
wire sgo__n315;
wire slo__n415;
wire sgo__n31;
wire sgo__n34;
wire sgo__n39;
wire slo___n553;
wire slo__n580;
wire sgo__n46;
wire sgo__n48;
wire sgo__n50;
wire slo__sro_n602;
wire drc_ipo_n910;
wire sgo__n66;
wire sgo__n69;
wire sgo__n74;
wire sgo__n106;
wire drc_ipo_n911;
wire sgo__n133;
wire sgo__n140;
wire sgo__n147;
wire sgo__n149;


AND2_X4 i_0_1098 (.ZN (\pp[0] [10] ), .A1 (y[10]), .A2 (x[0]));
BUF_X1 slo___L1_c736 (.Z (slo___n701), .A (n_0_4));
AND2_X4 i_0_1096 (.ZN (\pp[3] [10] ), .A1 (x[3]), .A2 (y[7]));
AND2_X4 i_0_1095 (.ZN (\pp[5] [10] ), .A1 (x[5]), .A2 (y[5]));
NAND2_X1 i_0_1094 (.ZN (n_0_74), .A1 (y[11]), .A2 (x[0]));
INV_X2 i_0_1093 (.ZN (\pp[0] [11] ), .A (n_0_74));
NAND2_X1 i_0_1092 (.ZN (n_0_73), .A1 (y[9]), .A2 (x[1]));
INV_X1 i_0_1091 (.ZN (\pp[1] [10] ), .A (n_0_73));
NAND2_X1 i_0_1090 (.ZN (n_0_72), .A1 (y[9]), .A2 (x[2]));
INV_X2 i_0_1089 (.ZN (\pp[2] [11] ), .A (n_0_72));
NAND2_X1 i_0_1088 (.ZN (n_0_71), .A1 (y[8]), .A2 (x[3]));
INV_X2 i_0_1067 (.ZN (\pp[3] [11] ), .A (n_0_71));
NAND2_X1 i_0_1066 (.ZN (n_0_70), .A1 (y[6]), .A2 (x[3]));
INV_X1 i_0_1055 (.ZN (\pp[3] [9] ), .A (n_0_70));
NAND2_X1 i_0_1032 (.ZN (n_0_69), .A1 (y[6]), .A2 (x[4]));
INV_X1 i_0_1022 (.ZN (\pp[4] [10] ), .A (n_0_69));
NAND2_X1 i_0_999 (.ZN (n_0_68), .A1 (y[6]), .A2 (x[5]));
INV_X2 i_0_998 (.ZN (\pp[5] [11] ), .A (n_0_68));
NAND2_X1 i_0_989 (.ZN (n_0_67), .A1 (y[4]), .A2 (x[5]));
INV_X2 i_0_965 (.ZN (\pp[5] [9] ), .A (n_0_67));
NAND2_X1 i_0_964 (.ZN (n_0_66), .A1 (y[4]), .A2 (x[6]));
INV_X2 i_0_963 (.ZN (\pp[6] [10] ), .A (n_0_66));
NAND2_X1 i_0_956 (.ZN (n_0_65), .A1 (y[3]), .A2 (x[6]));
INV_X1 i_0_930 (.ZN (\pp[6] [9] ), .A (n_0_65));
NAND2_X1 i_0_923 (.ZN (n_0_64), .A1 (y[2]), .A2 (x[8]));
INV_X1 i_0_897 (.ZN (\pp[8] [10] ), .A (n_0_64));
INV_X4 i_0_896 (.ZN (n_0_4), .A (y[2]));
INV_X16 i_0_895 (.ZN (n_0_5), .A (y[3]));
INV_X4 i_0_890 (.ZN (n_0_6), .A (y[4]));
INV_X16 i_0_862 (.ZN (n_0_7), .A (y[5]));
INV_X4 i_0_861 (.ZN (n_0_8), .A (y[6]));
INV_X4 i_0_857 (.ZN (n_0_9), .A (y[7]));
INV_X8 i_0_794 (.ZN (n_0_10), .A (y[8]));
INV_X4 i_0_791 (.ZN (n_0_11), .A (y[9]));
INV_X4 i_0_56 (.ZN (n_0_12), .A (y[10]));
INV_X8 i_0_54 (.ZN (n_0_13), .A (y[11]));
INV_X8 i_0_52 (.ZN (n_0_55), .A (x[8]));
INV_X8 i_0_50 (.ZN (n_0_57), .A (x[6]));
INV_X4 i_0_48 (.ZN (n_0_58), .A (x[5]));
INV_X8 i_0_46 (.ZN (n_0_59), .A (x[4]));
INV_X16 i_0_44 (.ZN (n_0_60), .A (x[3]));
INV_X8 i_0_42 (.ZN (n_0_61), .A (x[2]));
INV_X8 i_0_40 (.ZN (n_0_62), .A (x[1]));
INV_X4 i_0_38 (.ZN (n_0_63), .A (x[0]));
NOR2_X1 i_0_1087 (.ZN (\pp[0] [63] ), .A1 (n_0_33), .A2 (sgo__n301));
NOR2_X1 i_0_1086 (.ZN (\pp[0] [30] ), .A1 (n_0_32), .A2 (sgo__n301));
NOR2_X1 i_0_1085 (.ZN (\pp[0] [29] ), .A1 (n_0_31), .A2 (sgo__n301));
NOR2_X1 i_0_1084 (.ZN (\pp[0] [28] ), .A1 (n_0_30), .A2 (sgo__n301));
NOR2_X1 i_0_1083 (.ZN (\pp[0] [27] ), .A1 (n_0_29), .A2 (sgo__n301));
NOR2_X1 i_0_1082 (.ZN (\pp[0] [26] ), .A1 (n_0_28), .A2 (sgo__n301));
NOR2_X1 i_0_1081 (.ZN (\pp[0] [25] ), .A1 (n_0_27), .A2 (sgo__n301));
NOR2_X1 i_0_1080 (.ZN (\pp[0] [24] ), .A1 (n_0_26), .A2 (sgo__n301));
NOR2_X1 i_0_1079 (.ZN (\pp[0] [23] ), .A1 (n_0_25), .A2 (sgo__n301));
NOR2_X1 i_0_1078 (.ZN (\pp[0] [22] ), .A1 (n_0_24), .A2 (sgo__n301));
NOR2_X1 i_0_1077 (.ZN (\pp[0] [21] ), .A1 (n_0_23), .A2 (sgo__n301));
NOR2_X1 i_0_1076 (.ZN (\pp[0] [20] ), .A1 (n_0_22), .A2 (sgo__n301));
NOR2_X1 i_0_1075 (.ZN (\pp[0] [19] ), .A1 (n_0_21), .A2 (sgo__n301));
NOR2_X1 i_0_1074 (.ZN (\pp[0] [18] ), .A1 (n_0_20), .A2 (sgo__n301));
NOR2_X1 i_0_1073 (.ZN (\pp[0] [17] ), .A1 (n_0_19), .A2 (sgo__n301));
NOR2_X1 i_0_1072 (.ZN (\pp[0] [16] ), .A1 (n_0_18), .A2 (sgo__n301));
NOR2_X2 i_0_1071 (.ZN (\pp[0] [15] ), .A1 (n_0_17), .A2 (n_0_63));
NOR2_X1 i_0_1070 (.ZN (\pp[0] [14] ), .A1 (n_0_16), .A2 (sgo__n301));
NOR2_X4 i_0_1069 (.ZN (\pp[0] [13] ), .A1 (n_0_15), .A2 (n_0_63));
NOR2_X2 i_0_1068 (.ZN (\pp[0] [12] ), .A1 (n_0_14), .A2 (n_0_63));
NOR2_X4 i_0_1065 (.ZN (\pp[0] [9] ), .A1 (n_0_11), .A2 (n_0_63));
NOR2_X4 i_0_1064 (.ZN (\pp[0] [8] ), .A1 (n_0_10), .A2 (n_0_63));
NOR2_X2 i_0_1063 (.ZN (\pp[0] [7] ), .A1 (n_0_9), .A2 (n_0_63));
NOR2_X4 i_0_1062 (.ZN (\pp[0] [6] ), .A1 (sgo__n184), .A2 (sgo__n301));
NOR2_X4 i_0_1061 (.ZN (\pp[0] [5] ), .A1 (sgo__n172), .A2 (n_0_63));
NOR2_X2 i_0_1060 (.ZN (\pp[0] [4] ), .A1 (sgo__n205), .A2 (sgo__n301));
NOR2_X2 i_0_1059 (.ZN (\pp[0] [3] ), .A1 (n_0_5), .A2 (sgo__n301));
NOR2_X2 i_0_1058 (.ZN (\pp[0] [2] ), .A1 (n_0_4), .A2 (sgo__n301));
NOR2_X1 i_0_1057 (.ZN (\pp[0] [1] ), .A1 (n_0_3), .A2 (sgo__n301));
NOR2_X1 i_0_1056 (.ZN (\pp[0] [0] ), .A1 (n_0_2), .A2 (sgo__n301));
NOR2_X1 i_0_1054 (.ZN (\pp[1] [63] ), .A1 (n_0_62), .A2 (n_0_33));
NOR2_X1 i_0_1053 (.ZN (\pp[1] [31] ), .A1 (n_0_62), .A2 (n_0_32));
NOR2_X1 i_0_1052 (.ZN (\pp[1] [30] ), .A1 (n_0_62), .A2 (n_0_31));
NOR2_X1 i_0_1051 (.ZN (\pp[1] [29] ), .A1 (n_0_62), .A2 (n_0_30));
NOR2_X1 i_0_1050 (.ZN (\pp[1] [28] ), .A1 (n_0_62), .A2 (n_0_29));
NOR2_X1 i_0_1049 (.ZN (\pp[1] [27] ), .A1 (n_0_62), .A2 (n_0_28));
NOR2_X1 i_0_1048 (.ZN (\pp[1] [26] ), .A1 (n_0_62), .A2 (n_0_27));
NOR2_X1 i_0_1047 (.ZN (\pp[1] [25] ), .A1 (n_0_62), .A2 (n_0_26));
NOR2_X1 i_0_1046 (.ZN (\pp[1] [24] ), .A1 (n_0_62), .A2 (n_0_25));
NOR2_X1 i_0_1045 (.ZN (\pp[1] [23] ), .A1 (n_0_62), .A2 (n_0_24));
NOR2_X1 i_0_1044 (.ZN (\pp[1] [22] ), .A1 (n_0_62), .A2 (n_0_23));
NOR2_X1 i_0_1043 (.ZN (\pp[1] [21] ), .A1 (n_0_62), .A2 (n_0_22));
NOR2_X1 i_0_1042 (.ZN (\pp[1] [20] ), .A1 (n_0_62), .A2 (n_0_21));
NOR2_X1 i_0_1041 (.ZN (\pp[1] [19] ), .A1 (n_0_62), .A2 (n_0_20));
NOR2_X1 i_0_1040 (.ZN (\pp[1] [18] ), .A1 (n_0_62), .A2 (n_0_19));
NOR2_X1 i_0_1039 (.ZN (\pp[1] [17] ), .A1 (n_0_62), .A2 (n_0_18));
NOR2_X1 i_0_1038 (.ZN (\pp[1] [16] ), .A1 (n_0_62), .A2 (n_0_17));
NOR2_X1 i_0_1037 (.ZN (\pp[1] [15] ), .A1 (n_0_62), .A2 (n_0_16));
NOR2_X1 i_0_1036 (.ZN (\pp[1] [14] ), .A1 (n_0_62), .A2 (sgo__n46));
NOR2_X1 i_0_1035 (.ZN (\pp[1] [13] ), .A1 (n_0_62), .A2 (n_0_14));
NOR2_X2 i_0_1034 (.ZN (\pp[1] [12] ), .A1 (n_0_62), .A2 (n_0_13));
NOR2_X4 i_0_1033 (.ZN (\pp[1] [11] ), .A1 (n_0_62), .A2 (n_0_12));
NOR2_X4 i_0_1031 (.ZN (\pp[1] [9] ), .A1 (n_0_62), .A2 (n_0_10));
NOR2_X1 i_0_1030 (.ZN (\pp[1] [8] ), .A1 (n_0_62), .A2 (n_0_9));
NOR2_X1 i_0_1029 (.ZN (\pp[1] [7] ), .A1 (n_0_62), .A2 (n_0_8));
NOR2_X1 i_0_1028 (.ZN (\pp[1] [6] ), .A1 (n_0_62), .A2 (sgo__n172));
NOR2_X1 i_0_1027 (.ZN (\pp[1] [5] ), .A1 (n_0_62), .A2 (sgo__n205));
NOR2_X1 i_0_1026 (.ZN (\pp[1] [4] ), .A1 (n_0_62), .A2 (n_0_5));
NOR2_X1 i_0_1025 (.ZN (\pp[1] [3] ), .A1 (n_0_62), .A2 (sgo__n66));
NOR2_X1 i_0_1024 (.ZN (\pp[1] [2] ), .A1 (n_0_62), .A2 (sgo__n31));
NOR2_X1 i_0_1023 (.ZN (\pp[1] [1] ), .A1 (n_0_62), .A2 (sgo__n39));
NOR2_X1 i_0_1021 (.ZN (\pp[2] [63] ), .A1 (sgo__n167), .A2 (n_0_33));
NOR2_X1 i_0_1020 (.ZN (\pp[2] [32] ), .A1 (sgo__n167), .A2 (n_0_32));
NOR2_X1 i_0_1019 (.ZN (\pp[2] [31] ), .A1 (sgo__n167), .A2 (n_0_31));
NOR2_X1 i_0_1018 (.ZN (\pp[2] [30] ), .A1 (sgo__n167), .A2 (n_0_30));
NOR2_X1 i_0_1017 (.ZN (\pp[2] [29] ), .A1 (sgo__n167), .A2 (n_0_29));
NOR2_X1 i_0_1016 (.ZN (\pp[2] [28] ), .A1 (sgo__n167), .A2 (n_0_28));
NOR2_X1 i_0_1015 (.ZN (\pp[2] [27] ), .A1 (sgo__n167), .A2 (n_0_27));
NOR2_X1 i_0_1014 (.ZN (\pp[2] [26] ), .A1 (sgo__n167), .A2 (n_0_26));
NOR2_X1 i_0_1013 (.ZN (\pp[2] [25] ), .A1 (sgo__n167), .A2 (n_0_25));
NOR2_X1 i_0_1012 (.ZN (\pp[2] [24] ), .A1 (sgo__n167), .A2 (n_0_24));
NOR2_X1 i_0_1011 (.ZN (\pp[2] [23] ), .A1 (sgo__n167), .A2 (n_0_23));
NOR2_X1 i_0_1010 (.ZN (\pp[2] [22] ), .A1 (sgo__n167), .A2 (n_0_22));
NOR2_X1 i_0_1009 (.ZN (\pp[2] [21] ), .A1 (sgo__n167), .A2 (n_0_21));
NOR2_X1 i_0_1008 (.ZN (\pp[2] [20] ), .A1 (sgo__n167), .A2 (n_0_20));
NOR2_X1 i_0_1007 (.ZN (\pp[2] [19] ), .A1 (sgo__n167), .A2 (n_0_19));
NOR2_X1 i_0_1006 (.ZN (\pp[2] [18] ), .A1 (sgo__n167), .A2 (n_0_18));
NOR2_X2 i_0_1005 (.ZN (\pp[2] [17] ), .A1 (sgo__n167), .A2 (n_0_17));
NOR2_X1 i_0_1004 (.ZN (\pp[2] [16] ), .A1 (sgo__n167), .A2 (n_0_16));
NOR2_X2 i_0_1003 (.ZN (\pp[2] [15] ), .A1 (n_0_61), .A2 (sgo__n46));
NOR2_X1 i_0_1002 (.ZN (\pp[2] [14] ), .A1 (n_0_61), .A2 (n_0_14));
NOR2_X4 i_0_1001 (.ZN (\pp[2] [13] ), .A1 (slo__n415), .A2 (n_0_13));
NOR2_X4 i_0_1000 (.ZN (\pp[2] [12] ), .A1 (n_0_61), .A2 (n_0_12));
NOR2_X4 i_0_997 (.ZN (\pp[2] [9] ), .A1 (n_0_61), .A2 (n_0_9));
NOR2_X4 i_0_996 (.ZN (\pp[2] [8] ), .A1 (n_0_8), .A2 (n_0_61));
NOR2_X4 i_0_995 (.ZN (\pp[2] [7] ), .A1 (slo__n415), .A2 (n_0_7));
NOR2_X1 i_0_994 (.ZN (\pp[2] [6] ), .A1 (slo__n415), .A2 (sgo__n149));
NOR2_X1 i_0_993 (.ZN (\pp[2] [5] ), .A1 (sgo__n167), .A2 (n_0_5));
NOR2_X1 i_0_992 (.ZN (\pp[2] [4] ), .A1 (sgo__n167), .A2 (sgo__n66));
NOR2_X1 i_0_991 (.ZN (\pp[2] [3] ), .A1 (sgo__n167), .A2 (sgo__n31));
NOR2_X1 i_0_990 (.ZN (\pp[2] [2] ), .A1 (sgo__n167), .A2 (sgo__n39));
NOR2_X1 i_0_988 (.ZN (\pp[3] [63] ), .A1 (sgo__n150), .A2 (n_0_33));
NOR2_X1 i_0_987 (.ZN (\pp[3] [33] ), .A1 (sgo__n150), .A2 (n_0_32));
NOR2_X1 i_0_986 (.ZN (\pp[3] [32] ), .A1 (sgo__n150), .A2 (n_0_31));
NOR2_X1 i_0_985 (.ZN (\pp[3] [31] ), .A1 (sgo__n150), .A2 (n_0_30));
NOR2_X1 i_0_984 (.ZN (\pp[3] [30] ), .A1 (sgo__n150), .A2 (n_0_29));
NOR2_X1 i_0_983 (.ZN (\pp[3] [29] ), .A1 (sgo__n150), .A2 (n_0_28));
NOR2_X1 i_0_982 (.ZN (\pp[3] [28] ), .A1 (sgo__n150), .A2 (n_0_27));
NOR2_X1 i_0_981 (.ZN (\pp[3] [27] ), .A1 (sgo__n150), .A2 (n_0_26));
NOR2_X1 i_0_980 (.ZN (\pp[3] [26] ), .A1 (sgo__n150), .A2 (n_0_25));
NOR2_X1 i_0_979 (.ZN (\pp[3] [25] ), .A1 (sgo__n150), .A2 (n_0_24));
NOR2_X1 i_0_978 (.ZN (\pp[3] [24] ), .A1 (sgo__n150), .A2 (n_0_23));
NOR2_X1 i_0_977 (.ZN (\pp[3] [23] ), .A1 (sgo__n150), .A2 (n_0_22));
NOR2_X1 i_0_976 (.ZN (\pp[3] [22] ), .A1 (sgo__n150), .A2 (n_0_21));
NOR2_X1 i_0_975 (.ZN (\pp[3] [21] ), .A1 (sgo__n150), .A2 (n_0_20));
NOR2_X1 i_0_974 (.ZN (\pp[3] [20] ), .A1 (sgo__n150), .A2 (n_0_19));
NOR2_X1 i_0_973 (.ZN (\pp[3] [19] ), .A1 (sgo__n150), .A2 (n_0_18));
NOR2_X1 i_0_972 (.ZN (\pp[3] [18] ), .A1 (sgo__n150), .A2 (n_0_17));
NOR2_X1 i_0_971 (.ZN (\pp[3] [17] ), .A1 (sgo__n150), .A2 (n_0_16));
NOR2_X2 i_0_970 (.ZN (\pp[3] [16] ), .A1 (sgo__n150), .A2 (sgo__n46));
NOR2_X1 i_0_969 (.ZN (\pp[3] [15] ), .A1 (sgo__n150), .A2 (n_0_14));
NOR2_X1 i_0_968 (.ZN (\pp[3] [14] ), .A1 (sgo__n150), .A2 (n_0_13));
NOR2_X4 i_0_967 (.ZN (\pp[3] [13] ), .A1 (n_0_60), .A2 (n_0_12));
NOR2_X2 i_0_966 (.ZN (\pp[3] [12] ), .A1 (n_0_60), .A2 (n_0_11));
NOR2_X2 i_0_962 (.ZN (\pp[3] [8] ), .A1 (n_0_60), .A2 (n_0_7));
NOR2_X4 i_0_961 (.ZN (\pp[3] [7] ), .A1 (n_0_60), .A2 (sgo__n149));
NOR2_X1 i_0_960 (.ZN (\pp[3] [6] ), .A1 (sgo__n150), .A2 (n_0_5));
NOR2_X1 i_0_959 (.ZN (\pp[3] [5] ), .A1 (sgo__n150), .A2 (sgo__n66));
NOR2_X1 i_0_958 (.ZN (\pp[3] [4] ), .A1 (sgo__n150), .A2 (sgo__n31));
NOR2_X1 i_0_957 (.ZN (\pp[3] [3] ), .A1 (sgo__n150), .A2 (sgo__n39));
NOR2_X1 i_0_955 (.ZN (\pp[4] [63] ), .A1 (sgo__n315), .A2 (n_0_33));
NOR2_X1 i_0_954 (.ZN (\pp[4] [34] ), .A1 (sgo__n315), .A2 (n_0_32));
NOR2_X1 i_0_953 (.ZN (\pp[4] [33] ), .A1 (sgo__n315), .A2 (n_0_31));
NOR2_X1 i_0_952 (.ZN (\pp[4] [32] ), .A1 (sgo__n315), .A2 (n_0_30));
NOR2_X1 i_0_951 (.ZN (\pp[4] [31] ), .A1 (sgo__n315), .A2 (n_0_29));
NOR2_X1 i_0_950 (.ZN (\pp[4] [30] ), .A1 (sgo__n315), .A2 (n_0_28));
NOR2_X1 i_0_949 (.ZN (\pp[4] [29] ), .A1 (sgo__n315), .A2 (n_0_27));
NOR2_X1 i_0_948 (.ZN (\pp[4] [28] ), .A1 (sgo__n315), .A2 (n_0_26));
NOR2_X1 i_0_947 (.ZN (\pp[4] [27] ), .A1 (sgo__n315), .A2 (n_0_25));
NOR2_X1 i_0_946 (.ZN (\pp[4] [26] ), .A1 (sgo__n315), .A2 (n_0_24));
NOR2_X1 i_0_945 (.ZN (\pp[4] [25] ), .A1 (sgo__n315), .A2 (n_0_23));
NOR2_X1 i_0_944 (.ZN (\pp[4] [24] ), .A1 (sgo__n315), .A2 (n_0_22));
NOR2_X1 i_0_943 (.ZN (\pp[4] [23] ), .A1 (sgo__n315), .A2 (n_0_21));
NOR2_X1 i_0_942 (.ZN (\pp[4] [22] ), .A1 (sgo__n315), .A2 (n_0_20));
NOR2_X1 i_0_941 (.ZN (\pp[4] [21] ), .A1 (sgo__n315), .A2 (n_0_19));
NOR2_X1 i_0_940 (.ZN (\pp[4] [20] ), .A1 (sgo__n315), .A2 (n_0_18));
NOR2_X1 i_0_939 (.ZN (\pp[4] [19] ), .A1 (sgo__n315), .A2 (n_0_17));
NOR2_X1 i_0_938 (.ZN (\pp[4] [18] ), .A1 (sgo__n315), .A2 (n_0_16));
NOR2_X1 i_0_937 (.ZN (\pp[4] [17] ), .A1 (sgo__n315), .A2 (sgo__n46));
NOR2_X1 i_0_936 (.ZN (\pp[4] [16] ), .A1 (sgo__n315), .A2 (n_0_14));
NOR2_X1 i_0_935 (.ZN (\pp[4] [15] ), .A1 (sgo__n315), .A2 (n_0_13));
NOR2_X1 i_0_934 (.ZN (\pp[4] [14] ), .A1 (sgo__n315), .A2 (sgo__n157));
NOR2_X1 i_0_933 (.ZN (\pp[4] [13] ), .A1 (sgo__n315), .A2 (sgo__n177));
NOR2_X1 i_0_932 (.ZN (\pp[4] [12] ), .A1 (n_0_59), .A2 (n_0_10));
NOR2_X2 i_0_931 (.ZN (\pp[4] [11] ), .A1 (n_0_59), .A2 (n_0_9));
NOR2_X4 i_0_929 (.ZN (\pp[4] [9] ), .A1 (n_0_59), .A2 (n_0_7));
NOR2_X1 i_0_928 (.ZN (\pp[4] [8] ), .A1 (slo__n580), .A2 (n_0_59));
NOR2_X1 i_0_927 (.ZN (\pp[4] [7] ), .A1 (n_0_59), .A2 (n_0_5));
NOR2_X1 i_0_926 (.ZN (\pp[4] [6] ), .A1 (sgo__n315), .A2 (sgo__n66));
NOR2_X1 i_0_925 (.ZN (\pp[4] [5] ), .A1 (sgo__n315), .A2 (sgo__n31));
NOR2_X1 i_0_924 (.ZN (\pp[4] [4] ), .A1 (sgo__n315), .A2 (sgo__n39));
NOR2_X1 i_0_922 (.ZN (\pp[5] [63] ), .A1 (slo___n552), .A2 (n_0_33));
NOR2_X1 i_0_921 (.ZN (\pp[5] [35] ), .A1 (slo___n552), .A2 (n_0_32));
NOR2_X1 i_0_920 (.ZN (\pp[5] [34] ), .A1 (slo___n552), .A2 (n_0_31));
NOR2_X1 i_0_919 (.ZN (\pp[5] [33] ), .A1 (n_0_58), .A2 (n_0_30));
NOR2_X1 i_0_918 (.ZN (\pp[5] [32] ), .A1 (n_0_58), .A2 (n_0_29));
NOR2_X1 i_0_917 (.ZN (\pp[5] [31] ), .A1 (n_0_58), .A2 (n_0_28));
NOR2_X1 i_0_916 (.ZN (\pp[5] [30] ), .A1 (n_0_58), .A2 (n_0_27));
NOR2_X1 i_0_915 (.ZN (\pp[5] [29] ), .A1 (n_0_58), .A2 (n_0_26));
NOR2_X1 i_0_914 (.ZN (\pp[5] [28] ), .A1 (n_0_58), .A2 (n_0_25));
NOR2_X1 i_0_913 (.ZN (\pp[5] [27] ), .A1 (n_0_58), .A2 (n_0_24));
NOR2_X1 i_0_912 (.ZN (\pp[5] [26] ), .A1 (n_0_58), .A2 (n_0_23));
NOR2_X1 i_0_911 (.ZN (\pp[5] [25] ), .A1 (n_0_58), .A2 (n_0_22));
NOR2_X1 i_0_910 (.ZN (\pp[5] [24] ), .A1 (n_0_58), .A2 (n_0_21));
NOR2_X1 i_0_909 (.ZN (\pp[5] [23] ), .A1 (n_0_58), .A2 (n_0_20));
NOR2_X1 i_0_908 (.ZN (\pp[5] [22] ), .A1 (n_0_58), .A2 (n_0_19));
NOR2_X1 i_0_907 (.ZN (\pp[5] [21] ), .A1 (n_0_58), .A2 (n_0_18));
NOR2_X1 i_0_906 (.ZN (\pp[5] [20] ), .A1 (n_0_58), .A2 (n_0_17));
NOR2_X1 i_0_905 (.ZN (\pp[5] [19] ), .A1 (n_0_58), .A2 (n_0_16));
NOR2_X1 i_0_904 (.ZN (\pp[5] [18] ), .A1 (n_0_58), .A2 (n_0_15));
NOR2_X1 i_0_903 (.ZN (\pp[5] [17] ), .A1 (n_0_58), .A2 (n_0_14));
NOR2_X1 i_0_902 (.ZN (\pp[5] [16] ), .A1 (n_0_58), .A2 (n_0_13));
NOR2_X4 i_0_901 (.ZN (\pp[5] [15] ), .A1 (n_0_58), .A2 (n_0_12));
NOR2_X1 i_0_900 (.ZN (\pp[5] [14] ), .A1 (n_0_58), .A2 (n_0_11));
NOR2_X2 i_0_899 (.ZN (\pp[5] [13] ), .A1 (n_0_58), .A2 (n_0_10));
NOR2_X4 i_0_898 (.ZN (\pp[5] [12] ), .A1 (n_0_58), .A2 (n_0_9));
NOR2_X2 i_0_894 (.ZN (\pp[5] [8] ), .A1 (n_0_58), .A2 (n_0_5));
NOR2_X2 i_0_893 (.ZN (\pp[5] [7] ), .A1 (n_0_58), .A2 (n_0_4));
NOR2_X2 i_0_892 (.ZN (\pp[5] [6] ), .A1 (slo___n553), .A2 (sgo__n31));
NOR2_X1 i_0_891 (.ZN (\pp[5] [5] ), .A1 (slo___n553), .A2 (sgo__n39));
NOR2_X1 i_0_889 (.ZN (\pp[6] [63] ), .A1 (n_0_57), .A2 (n_0_33));
NOR2_X1 i_0_888 (.ZN (\pp[6] [36] ), .A1 (n_0_57), .A2 (n_0_32));
NOR2_X1 i_0_887 (.ZN (\pp[6] [35] ), .A1 (n_0_57), .A2 (n_0_31));
NOR2_X1 i_0_886 (.ZN (\pp[6] [34] ), .A1 (n_0_57), .A2 (n_0_30));
NOR2_X1 i_0_885 (.ZN (\pp[6] [33] ), .A1 (n_0_57), .A2 (n_0_29));
NOR2_X1 i_0_884 (.ZN (\pp[6] [32] ), .A1 (n_0_57), .A2 (n_0_28));
NOR2_X1 i_0_883 (.ZN (\pp[6] [31] ), .A1 (n_0_57), .A2 (n_0_27));
NOR2_X1 i_0_882 (.ZN (\pp[6] [30] ), .A1 (n_0_57), .A2 (n_0_26));
NOR2_X1 i_0_881 (.ZN (\pp[6] [29] ), .A1 (n_0_57), .A2 (n_0_25));
NOR2_X1 i_0_880 (.ZN (\pp[6] [28] ), .A1 (n_0_57), .A2 (n_0_24));
NOR2_X1 i_0_879 (.ZN (\pp[6] [27] ), .A1 (n_0_57), .A2 (n_0_23));
NOR2_X1 i_0_878 (.ZN (\pp[6] [26] ), .A1 (n_0_57), .A2 (n_0_22));
NOR2_X1 i_0_877 (.ZN (\pp[6] [25] ), .A1 (n_0_57), .A2 (n_0_21));
NOR2_X1 i_0_876 (.ZN (\pp[6] [24] ), .A1 (n_0_57), .A2 (n_0_20));
NOR2_X1 i_0_875 (.ZN (\pp[6] [23] ), .A1 (n_0_57), .A2 (n_0_19));
NOR2_X1 i_0_874 (.ZN (\pp[6] [22] ), .A1 (n_0_57), .A2 (n_0_18));
NOR2_X1 i_0_873 (.ZN (\pp[6] [21] ), .A1 (n_0_57), .A2 (n_0_17));
NOR2_X1 i_0_872 (.ZN (\pp[6] [20] ), .A1 (n_0_57), .A2 (n_0_16));
NOR2_X1 i_0_871 (.ZN (\pp[6] [19] ), .A1 (n_0_57), .A2 (sgo__n48));
NOR2_X1 i_0_870 (.ZN (\pp[6] [18] ), .A1 (n_0_57), .A2 (sgo__n240));
NOR2_X1 i_0_869 (.ZN (\pp[6] [17] ), .A1 (n_0_57), .A2 (n_0_13));
NOR2_X1 i_0_868 (.ZN (\pp[6] [16] ), .A1 (n_0_57), .A2 (sgo__n157));
NOR2_X1 i_0_867 (.ZN (\pp[6] [15] ), .A1 (n_0_57), .A2 (sgo__n177));
NOR2_X1 i_0_866 (.ZN (\pp[6] [14] ), .A1 (n_0_57), .A2 (sgo__n162));
NOR2_X1 i_0_865 (.ZN (\pp[6] [13] ), .A1 (n_0_57), .A2 (n_0_9));
NOR2_X2 i_0_864 (.ZN (\pp[6] [12] ), .A1 (n_0_57), .A2 (n_0_8));
NOR2_X4 i_0_863 (.ZN (\pp[6] [11] ), .A1 (n_0_57), .A2 (n_0_7));
NOR2_X2 i_0_860 (.ZN (\pp[6] [8] ), .A1 (n_0_57), .A2 (n_0_4));
NOR2_X1 i_0_859 (.ZN (\pp[6] [7] ), .A1 (n_0_57), .A2 (n_0_3));
NOR2_X1 i_0_858 (.ZN (\pp[6] [6] ), .A1 (n_0_57), .A2 (sgo__n39));
NOR2_X1 i_0_856 (.ZN (\pp[7] [63] ), .A1 (n_0_56), .A2 (n_0_33));
NOR2_X1 i_0_855 (.ZN (\pp[7] [37] ), .A1 (n_0_56), .A2 (n_0_32));
NOR2_X1 i_0_854 (.ZN (\pp[7] [36] ), .A1 (n_0_56), .A2 (n_0_31));
NOR2_X1 i_0_853 (.ZN (\pp[7] [35] ), .A1 (n_0_56), .A2 (n_0_30));
NOR2_X1 i_0_852 (.ZN (\pp[7] [34] ), .A1 (n_0_56), .A2 (n_0_29));
NOR2_X1 i_0_851 (.ZN (\pp[7] [33] ), .A1 (n_0_56), .A2 (n_0_28));
NOR2_X1 i_0_850 (.ZN (\pp[7] [32] ), .A1 (n_0_56), .A2 (n_0_27));
NOR2_X1 i_0_849 (.ZN (\pp[7] [31] ), .A1 (n_0_56), .A2 (n_0_26));
NOR2_X1 i_0_848 (.ZN (\pp[7] [30] ), .A1 (n_0_56), .A2 (n_0_25));
NOR2_X1 i_0_847 (.ZN (\pp[7] [29] ), .A1 (n_0_56), .A2 (n_0_24));
NOR2_X1 i_0_846 (.ZN (\pp[7] [28] ), .A1 (n_0_56), .A2 (n_0_23));
NOR2_X1 i_0_845 (.ZN (\pp[7] [27] ), .A1 (n_0_56), .A2 (n_0_22));
NOR2_X1 i_0_844 (.ZN (\pp[7] [26] ), .A1 (n_0_56), .A2 (n_0_21));
NOR2_X1 i_0_843 (.ZN (\pp[7] [25] ), .A1 (n_0_56), .A2 (n_0_20));
NOR2_X1 i_0_842 (.ZN (\pp[7] [24] ), .A1 (n_0_56), .A2 (n_0_19));
NOR2_X1 i_0_841 (.ZN (\pp[7] [23] ), .A1 (n_0_56), .A2 (n_0_18));
NOR2_X1 i_0_840 (.ZN (\pp[7] [22] ), .A1 (n_0_56), .A2 (n_0_17));
NOR2_X1 i_0_839 (.ZN (\pp[7] [21] ), .A1 (n_0_56), .A2 (n_0_16));
NOR2_X1 i_0_838 (.ZN (\pp[7] [20] ), .A1 (n_0_56), .A2 (sgo__n48));
NOR2_X1 i_0_837 (.ZN (\pp[7] [19] ), .A1 (n_0_56), .A2 (sgo__n240));
NOR2_X1 i_0_836 (.ZN (\pp[7] [18] ), .A1 (n_0_56), .A2 (n_0_13));
NOR2_X1 i_0_835 (.ZN (\pp[7] [17] ), .A1 (n_0_56), .A2 (sgo__n157));
NOR2_X1 i_0_834 (.ZN (\pp[7] [16] ), .A1 (n_0_56), .A2 (sgo__n177));
NOR2_X1 i_0_833 (.ZN (\pp[7] [15] ), .A1 (n_0_56), .A2 (sgo__n162));
NOR2_X4 i_0_832 (.ZN (\pp[7] [14] ), .A1 (n_0_56), .A2 (n_0_9));
NOR2_X2 i_0_831 (.ZN (\pp[7] [13] ), .A1 (n_0_56), .A2 (sgo__n184));
NOR2_X2 i_0_830 (.ZN (\pp[7] [12] ), .A1 (n_0_56), .A2 (sgo__n172));
NOR2_X2 i_0_829 (.ZN (\pp[7] [11] ), .A1 (n_0_56), .A2 (n_0_6));
NOR2_X2 i_0_828 (.ZN (\pp[7] [10] ), .A1 (n_0_56), .A2 (n_0_5));
NOR2_X4 i_0_827 (.ZN (\pp[7] [9] ), .A1 (n_0_4), .A2 (n_0_56));
NOR2_X1 i_0_826 (.ZN (\pp[7] [8] ), .A1 (n_0_56), .A2 (n_0_3));
NOR2_X1 i_0_825 (.ZN (\pp[7] [7] ), .A1 (n_0_56), .A2 (n_0_2));
INV_X16 i_0_824 (.ZN (n_0_56), .A (x[7]));
NOR2_X1 i_0_823 (.ZN (\pp[8] [63] ), .A1 (sgo__n272), .A2 (n_0_33));
NOR2_X1 i_0_822 (.ZN (\pp[8] [38] ), .A1 (sgo__n272), .A2 (n_0_32));
NOR2_X1 i_0_821 (.ZN (\pp[8] [37] ), .A1 (sgo__n272), .A2 (n_0_31));
NOR2_X1 i_0_820 (.ZN (\pp[8] [36] ), .A1 (sgo__n272), .A2 (n_0_30));
NOR2_X1 i_0_819 (.ZN (\pp[8] [35] ), .A1 (sgo__n272), .A2 (n_0_29));
NOR2_X1 i_0_818 (.ZN (\pp[8] [34] ), .A1 (sgo__n272), .A2 (n_0_28));
NOR2_X1 i_0_817 (.ZN (\pp[8] [33] ), .A1 (sgo__n272), .A2 (n_0_27));
NOR2_X1 i_0_816 (.ZN (\pp[8] [32] ), .A1 (sgo__n272), .A2 (n_0_26));
NOR2_X1 i_0_815 (.ZN (\pp[8] [31] ), .A1 (sgo__n272), .A2 (n_0_25));
NOR2_X1 i_0_814 (.ZN (\pp[8] [30] ), .A1 (sgo__n272), .A2 (n_0_24));
NOR2_X1 i_0_813 (.ZN (\pp[8] [29] ), .A1 (sgo__n272), .A2 (n_0_23));
NOR2_X1 i_0_812 (.ZN (\pp[8] [28] ), .A1 (sgo__n272), .A2 (n_0_22));
NOR2_X1 i_0_811 (.ZN (\pp[8] [27] ), .A1 (sgo__n272), .A2 (n_0_21));
NOR2_X1 i_0_810 (.ZN (\pp[8] [26] ), .A1 (sgo__n272), .A2 (n_0_20));
NOR2_X1 i_0_809 (.ZN (\pp[8] [25] ), .A1 (sgo__n272), .A2 (n_0_19));
NOR2_X1 i_0_808 (.ZN (\pp[8] [24] ), .A1 (sgo__n272), .A2 (n_0_18));
NOR2_X1 i_0_807 (.ZN (\pp[8] [23] ), .A1 (sgo__n272), .A2 (n_0_17));
NOR2_X1 i_0_806 (.ZN (\pp[8] [22] ), .A1 (sgo__n272), .A2 (n_0_16));
NOR2_X1 i_0_805 (.ZN (\pp[8] [21] ), .A1 (sgo__n272), .A2 (sgo__n48));
NOR2_X1 i_0_804 (.ZN (\pp[8] [20] ), .A1 (sgo__n272), .A2 (sgo__n240));
NOR2_X1 i_0_803 (.ZN (\pp[8] [19] ), .A1 (sgo__n272), .A2 (n_0_13));
NOR2_X1 i_0_802 (.ZN (\pp[8] [18] ), .A1 (sgo__n272), .A2 (sgo__n157));
NOR2_X1 i_0_801 (.ZN (\pp[8] [17] ), .A1 (sgo__n272), .A2 (sgo__n177));
NOR2_X1 i_0_800 (.ZN (\pp[8] [16] ), .A1 (sgo__n272), .A2 (sgo__n162));
NOR2_X1 i_0_799 (.ZN (\pp[8] [15] ), .A1 (sgo__n272), .A2 (n_0_9));
NOR2_X2 i_0_798 (.ZN (\pp[8] [14] ), .A1 (sgo__n272), .A2 (sgo__n184));
NOR2_X2 i_0_797 (.ZN (\pp[8] [13] ), .A1 (sgo__n272), .A2 (sgo__n172));
NOR2_X2 i_0_796 (.ZN (\pp[8] [12] ), .A1 (n_0_55), .A2 (n_0_6));
NOR2_X2 i_0_795 (.ZN (\pp[8] [11] ), .A1 (n_0_55), .A2 (n_0_5));
NOR2_X4 i_0_793 (.ZN (\pp[8] [9] ), .A1 (n_0_3), .A2 (n_0_55));
NOR2_X4 i_0_792 (.ZN (\pp[8] [8] ), .A1 (n_0_55), .A2 (n_0_2));
NOR2_X1 i_0_790 (.ZN (\pp[9] [63] ), .A1 (n_0_54), .A2 (n_0_33));
NOR2_X1 i_0_789 (.ZN (\pp[9] [39] ), .A1 (n_0_54), .A2 (n_0_32));
NOR2_X1 i_0_788 (.ZN (\pp[9] [38] ), .A1 (n_0_54), .A2 (n_0_31));
NOR2_X1 i_0_787 (.ZN (\pp[9] [37] ), .A1 (n_0_54), .A2 (n_0_30));
NOR2_X1 i_0_786 (.ZN (\pp[9] [36] ), .A1 (n_0_54), .A2 (n_0_29));
NOR2_X1 i_0_785 (.ZN (\pp[9] [35] ), .A1 (n_0_54), .A2 (n_0_28));
NOR2_X1 i_0_784 (.ZN (\pp[9] [34] ), .A1 (n_0_54), .A2 (n_0_27));
NOR2_X1 i_0_783 (.ZN (\pp[9] [33] ), .A1 (n_0_54), .A2 (n_0_26));
NOR2_X1 i_0_782 (.ZN (\pp[9] [32] ), .A1 (n_0_54), .A2 (n_0_25));
NOR2_X1 i_0_781 (.ZN (\pp[9] [31] ), .A1 (n_0_54), .A2 (n_0_24));
NOR2_X1 i_0_780 (.ZN (\pp[9] [30] ), .A1 (n_0_54), .A2 (n_0_23));
NOR2_X1 i_0_779 (.ZN (\pp[9] [29] ), .A1 (n_0_54), .A2 (n_0_22));
NOR2_X1 i_0_778 (.ZN (\pp[9] [28] ), .A1 (n_0_54), .A2 (n_0_21));
NOR2_X1 i_0_777 (.ZN (\pp[9] [27] ), .A1 (n_0_54), .A2 (n_0_20));
NOR2_X1 i_0_776 (.ZN (\pp[9] [26] ), .A1 (n_0_54), .A2 (n_0_19));
NOR2_X1 i_0_775 (.ZN (\pp[9] [25] ), .A1 (n_0_54), .A2 (n_0_18));
NOR2_X1 i_0_774 (.ZN (\pp[9] [24] ), .A1 (n_0_54), .A2 (n_0_17));
NOR2_X1 i_0_773 (.ZN (\pp[9] [23] ), .A1 (n_0_54), .A2 (n_0_16));
NOR2_X1 i_0_772 (.ZN (\pp[9] [22] ), .A1 (n_0_54), .A2 (n_0_15));
NOR2_X1 i_0_771 (.ZN (\pp[9] [21] ), .A1 (n_0_54), .A2 (sgo__n240));
NOR2_X1 i_0_770 (.ZN (\pp[9] [20] ), .A1 (n_0_54), .A2 (n_0_13));
NOR2_X1 i_0_769 (.ZN (\pp[9] [19] ), .A1 (n_0_54), .A2 (sgo__n157));
NOR2_X1 i_0_768 (.ZN (\pp[9] [18] ), .A1 (n_0_54), .A2 (sgo__n177));
NOR2_X1 i_0_767 (.ZN (\pp[9] [17] ), .A1 (n_0_54), .A2 (sgo__n162));
NOR2_X1 i_0_766 (.ZN (\pp[9] [16] ), .A1 (n_0_54), .A2 (n_0_9));
NOR2_X2 i_0_765 (.ZN (\pp[9] [15] ), .A1 (n_0_54), .A2 (sgo__n184));
NOR2_X2 i_0_764 (.ZN (\pp[9] [14] ), .A1 (n_0_54), .A2 (sgo__n172));
NOR2_X2 i_0_763 (.ZN (\pp[9] [13] ), .A1 (n_0_54), .A2 (sgo__n149));
NOR2_X2 i_0_762 (.ZN (\pp[9] [12] ), .A1 (n_0_54), .A2 (n_0_5));
BUF_X1 slo___L1_c590 (.Z (slo___n552), .A (n_0_58));
NOR2_X1 i_0_760 (.ZN (\pp[9] [10] ), .A1 (n_0_54), .A2 (n_0_3));
NOR2_X1 i_0_759 (.ZN (\pp[9] [9] ), .A1 (n_0_54), .A2 (n_0_2));
INV_X8 i_0_758 (.ZN (n_0_54), .A (x[9]));
NOR2_X1 i_0_757 (.ZN (\pp[10] [63] ), .A1 (n_0_53), .A2 (n_0_33));
NOR2_X1 i_0_756 (.ZN (\pp[10] [40] ), .A1 (n_0_53), .A2 (n_0_32));
NOR2_X1 i_0_755 (.ZN (\pp[10] [39] ), .A1 (n_0_53), .A2 (n_0_31));
NOR2_X1 i_0_754 (.ZN (\pp[10] [38] ), .A1 (n_0_53), .A2 (n_0_30));
NOR2_X1 i_0_753 (.ZN (\pp[10] [37] ), .A1 (n_0_53), .A2 (n_0_29));
NOR2_X1 i_0_752 (.ZN (\pp[10] [36] ), .A1 (n_0_53), .A2 (n_0_28));
NOR2_X1 i_0_751 (.ZN (\pp[10] [35] ), .A1 (n_0_53), .A2 (n_0_27));
NOR2_X1 i_0_750 (.ZN (\pp[10] [34] ), .A1 (n_0_53), .A2 (n_0_26));
NOR2_X1 i_0_749 (.ZN (\pp[10] [33] ), .A1 (n_0_53), .A2 (n_0_25));
NOR2_X1 i_0_748 (.ZN (\pp[10] [32] ), .A1 (n_0_53), .A2 (n_0_24));
NOR2_X1 i_0_747 (.ZN (\pp[10] [31] ), .A1 (n_0_53), .A2 (n_0_23));
NOR2_X1 i_0_746 (.ZN (\pp[10] [30] ), .A1 (n_0_53), .A2 (n_0_22));
NOR2_X1 i_0_745 (.ZN (\pp[10] [29] ), .A1 (n_0_53), .A2 (n_0_21));
NOR2_X1 i_0_744 (.ZN (\pp[10] [28] ), .A1 (n_0_53), .A2 (n_0_20));
NOR2_X1 i_0_743 (.ZN (\pp[10] [27] ), .A1 (n_0_53), .A2 (n_0_19));
NOR2_X1 i_0_742 (.ZN (\pp[10] [26] ), .A1 (n_0_53), .A2 (n_0_18));
NOR2_X1 i_0_741 (.ZN (\pp[10] [25] ), .A1 (n_0_53), .A2 (n_0_17));
NOR2_X1 i_0_740 (.ZN (\pp[10] [24] ), .A1 (n_0_53), .A2 (n_0_16));
NOR2_X1 i_0_739 (.ZN (\pp[10] [23] ), .A1 (n_0_53), .A2 (n_0_15));
NOR2_X1 i_0_738 (.ZN (\pp[10] [22] ), .A1 (n_0_53), .A2 (sgo__n240));
NOR2_X1 i_0_737 (.ZN (\pp[10] [21] ), .A1 (n_0_53), .A2 (n_0_13));
NOR2_X1 i_0_736 (.ZN (\pp[10] [20] ), .A1 (n_0_53), .A2 (sgo__n157));
NOR2_X1 i_0_735 (.ZN (\pp[10] [19] ), .A1 (n_0_53), .A2 (sgo__n177));
NOR2_X1 i_0_734 (.ZN (\pp[10] [18] ), .A1 (n_0_53), .A2 (sgo__n162));
NOR2_X1 i_0_733 (.ZN (\pp[10] [17] ), .A1 (n_0_53), .A2 (n_0_9));
NOR2_X1 i_0_732 (.ZN (\pp[10] [16] ), .A1 (n_0_53), .A2 (sgo__n184));
NOR2_X1 i_0_731 (.ZN (\pp[10] [15] ), .A1 (n_0_53), .A2 (sgo__n172));
NOR2_X1 i_0_730 (.ZN (\pp[10] [14] ), .A1 (n_0_53), .A2 (sgo__n205));
NOR2_X1 i_0_729 (.ZN (\pp[10] [13] ), .A1 (n_0_53), .A2 (n_0_5));
NOR2_X1 i_0_728 (.ZN (\pp[10] [12] ), .A1 (n_0_53), .A2 (sgo__n66));
NOR2_X1 i_0_727 (.ZN (\pp[10] [11] ), .A1 (n_0_53), .A2 (n_0_3));
NOR2_X1 i_0_726 (.ZN (\pp[10] [10] ), .A1 (n_0_53), .A2 (n_0_2));
INV_X16 i_0_725 (.ZN (n_0_53), .A (x[10]));
NOR2_X1 i_0_724 (.ZN (\pp[11] [63] ), .A1 (n_0_52), .A2 (n_0_33));
NOR2_X1 i_0_723 (.ZN (\pp[11] [41] ), .A1 (n_0_52), .A2 (n_0_32));
NOR2_X1 i_0_722 (.ZN (\pp[11] [40] ), .A1 (n_0_52), .A2 (n_0_31));
NOR2_X1 i_0_721 (.ZN (\pp[11] [39] ), .A1 (n_0_52), .A2 (n_0_30));
NOR2_X1 i_0_720 (.ZN (\pp[11] [38] ), .A1 (n_0_52), .A2 (n_0_29));
NOR2_X1 i_0_719 (.ZN (\pp[11] [37] ), .A1 (n_0_52), .A2 (n_0_28));
NOR2_X1 i_0_718 (.ZN (\pp[11] [36] ), .A1 (n_0_52), .A2 (n_0_27));
NOR2_X1 i_0_717 (.ZN (\pp[11] [35] ), .A1 (n_0_52), .A2 (n_0_26));
NOR2_X1 i_0_716 (.ZN (\pp[11] [34] ), .A1 (n_0_52), .A2 (n_0_25));
NOR2_X1 i_0_715 (.ZN (\pp[11] [33] ), .A1 (n_0_52), .A2 (n_0_24));
NOR2_X1 i_0_714 (.ZN (\pp[11] [32] ), .A1 (n_0_52), .A2 (n_0_23));
NOR2_X1 i_0_713 (.ZN (\pp[11] [31] ), .A1 (n_0_52), .A2 (n_0_22));
NOR2_X1 i_0_712 (.ZN (\pp[11] [30] ), .A1 (n_0_52), .A2 (n_0_21));
NOR2_X1 i_0_711 (.ZN (\pp[11] [29] ), .A1 (n_0_52), .A2 (n_0_20));
NOR2_X1 i_0_710 (.ZN (\pp[11] [28] ), .A1 (n_0_52), .A2 (n_0_19));
NOR2_X1 i_0_709 (.ZN (\pp[11] [27] ), .A1 (n_0_52), .A2 (n_0_18));
NOR2_X1 i_0_708 (.ZN (\pp[11] [26] ), .A1 (n_0_52), .A2 (n_0_17));
NOR2_X1 i_0_707 (.ZN (\pp[11] [25] ), .A1 (n_0_52), .A2 (n_0_16));
NOR2_X1 i_0_706 (.ZN (\pp[11] [24] ), .A1 (n_0_52), .A2 (n_0_15));
NOR2_X1 i_0_705 (.ZN (\pp[11] [23] ), .A1 (n_0_52), .A2 (sgo__n240));
NOR2_X1 i_0_704 (.ZN (\pp[11] [22] ), .A1 (n_0_52), .A2 (n_0_13));
NOR2_X1 i_0_703 (.ZN (\pp[11] [21] ), .A1 (n_0_52), .A2 (sgo__n157));
NOR2_X1 i_0_702 (.ZN (\pp[11] [20] ), .A1 (n_0_52), .A2 (sgo__n177));
NOR2_X1 i_0_701 (.ZN (\pp[11] [19] ), .A1 (n_0_52), .A2 (sgo__n162));
NOR2_X1 i_0_700 (.ZN (\pp[11] [18] ), .A1 (n_0_52), .A2 (n_0_9));
NOR2_X1 i_0_699 (.ZN (\pp[11] [17] ), .A1 (n_0_52), .A2 (sgo__n184));
NOR2_X1 i_0_698 (.ZN (\pp[11] [16] ), .A1 (n_0_52), .A2 (sgo__n172));
NOR2_X2 i_0_697 (.ZN (\pp[11] [15] ), .A1 (n_0_52), .A2 (sgo__n205));
NOR2_X1 i_0_696 (.ZN (\pp[11] [14] ), .A1 (n_0_52), .A2 (n_0_5));
NOR2_X2 i_0_695 (.ZN (\pp[11] [13] ), .A1 (n_0_52), .A2 (sgo__n66));
NOR2_X4 i_0_693 (.ZN (\pp[11] [11] ), .A1 (n_0_52), .A2 (n_0_2));
INV_X16 i_0_692 (.ZN (n_0_52), .A (x[11]));
NOR2_X1 i_0_691 (.ZN (\pp[12] [62] ), .A1 (n_0_51), .A2 (n_0_33));
NOR2_X1 i_0_690 (.ZN (\pp[12] [42] ), .A1 (n_0_51), .A2 (n_0_32));
NOR2_X1 i_0_689 (.ZN (\pp[12] [41] ), .A1 (n_0_51), .A2 (n_0_31));
NOR2_X1 i_0_688 (.ZN (\pp[12] [40] ), .A1 (n_0_51), .A2 (n_0_30));
NOR2_X1 i_0_687 (.ZN (\pp[12] [39] ), .A1 (n_0_51), .A2 (n_0_29));
NOR2_X1 i_0_686 (.ZN (\pp[12] [38] ), .A1 (n_0_51), .A2 (n_0_28));
NOR2_X1 i_0_685 (.ZN (\pp[12] [37] ), .A1 (n_0_51), .A2 (n_0_27));
NOR2_X1 i_0_684 (.ZN (\pp[12] [36] ), .A1 (n_0_51), .A2 (n_0_26));
NOR2_X1 i_0_683 (.ZN (\pp[12] [35] ), .A1 (n_0_51), .A2 (n_0_25));
NOR2_X1 i_0_682 (.ZN (\pp[12] [34] ), .A1 (n_0_51), .A2 (n_0_24));
NOR2_X1 i_0_681 (.ZN (\pp[12] [33] ), .A1 (n_0_51), .A2 (n_0_23));
NOR2_X1 i_0_680 (.ZN (\pp[12] [32] ), .A1 (n_0_51), .A2 (n_0_22));
NOR2_X1 i_0_679 (.ZN (\pp[12] [31] ), .A1 (n_0_51), .A2 (n_0_21));
NOR2_X1 i_0_678 (.ZN (\pp[12] [30] ), .A1 (n_0_51), .A2 (n_0_20));
NOR2_X1 i_0_677 (.ZN (\pp[12] [29] ), .A1 (n_0_51), .A2 (n_0_19));
NOR2_X1 i_0_676 (.ZN (\pp[12] [28] ), .A1 (n_0_51), .A2 (n_0_18));
NOR2_X1 i_0_675 (.ZN (\pp[12] [27] ), .A1 (n_0_51), .A2 (n_0_17));
NOR2_X1 i_0_674 (.ZN (\pp[12] [26] ), .A1 (n_0_51), .A2 (n_0_16));
NOR2_X1 i_0_673 (.ZN (\pp[12] [25] ), .A1 (n_0_51), .A2 (n_0_15));
NOR2_X1 i_0_672 (.ZN (\pp[12] [24] ), .A1 (n_0_51), .A2 (sgo__n240));
NOR2_X1 i_0_671 (.ZN (\pp[12] [23] ), .A1 (n_0_51), .A2 (n_0_13));
NOR2_X1 i_0_670 (.ZN (\pp[12] [22] ), .A1 (n_0_51), .A2 (sgo__n157));
NOR2_X1 i_0_669 (.ZN (\pp[12] [21] ), .A1 (n_0_51), .A2 (sgo__n177));
NOR2_X1 i_0_668 (.ZN (\pp[12] [20] ), .A1 (n_0_51), .A2 (sgo__n162));
NOR2_X1 i_0_667 (.ZN (\pp[12] [19] ), .A1 (n_0_51), .A2 (n_0_9));
NOR2_X1 i_0_666 (.ZN (\pp[12] [18] ), .A1 (n_0_51), .A2 (sgo__n184));
NOR2_X1 i_0_665 (.ZN (\pp[12] [17] ), .A1 (n_0_51), .A2 (sgo__n172));
NOR2_X1 i_0_664 (.ZN (\pp[12] [16] ), .A1 (n_0_51), .A2 (sgo__n205));
NOR2_X2 i_0_663 (.ZN (\pp[12] [15] ), .A1 (n_0_51), .A2 (n_0_5));
NOR2_X2 i_0_662 (.ZN (\pp[12] [14] ), .A1 (n_0_51), .A2 (sgo__n66));
NOR2_X1 i_0_661 (.ZN (\pp[12] [13] ), .A1 (n_0_51), .A2 (sgo__n31));
NOR2_X1 i_0_660 (.ZN (\pp[12] [12] ), .A1 (n_0_51), .A2 (sgo__n39));
INV_X16 i_0_659 (.ZN (n_0_51), .A (x[12]));
NOR2_X1 i_0_658 (.ZN (\pp[13] [62] ), .A1 (n_0_50), .A2 (n_0_33));
NOR2_X1 i_0_657 (.ZN (\pp[13] [43] ), .A1 (n_0_50), .A2 (n_0_32));
NOR2_X1 i_0_656 (.ZN (\pp[13] [42] ), .A1 (n_0_50), .A2 (n_0_31));
NOR2_X1 i_0_655 (.ZN (\pp[13] [41] ), .A1 (n_0_50), .A2 (n_0_30));
NOR2_X1 i_0_654 (.ZN (\pp[13] [40] ), .A1 (n_0_50), .A2 (n_0_29));
NOR2_X1 i_0_653 (.ZN (\pp[13] [39] ), .A1 (n_0_50), .A2 (n_0_28));
NOR2_X1 i_0_652 (.ZN (\pp[13] [38] ), .A1 (n_0_50), .A2 (n_0_27));
NOR2_X1 i_0_651 (.ZN (\pp[13] [37] ), .A1 (n_0_50), .A2 (n_0_26));
NOR2_X1 i_0_650 (.ZN (\pp[13] [36] ), .A1 (n_0_50), .A2 (n_0_25));
NOR2_X1 i_0_649 (.ZN (\pp[13] [35] ), .A1 (n_0_50), .A2 (n_0_24));
NOR2_X1 i_0_648 (.ZN (\pp[13] [34] ), .A1 (n_0_50), .A2 (n_0_23));
NOR2_X1 i_0_647 (.ZN (\pp[13] [33] ), .A1 (n_0_50), .A2 (n_0_22));
NOR2_X1 i_0_646 (.ZN (\pp[13] [32] ), .A1 (n_0_50), .A2 (n_0_21));
NOR2_X1 i_0_645 (.ZN (\pp[13] [31] ), .A1 (n_0_50), .A2 (n_0_20));
NOR2_X1 i_0_644 (.ZN (\pp[13] [30] ), .A1 (n_0_50), .A2 (n_0_19));
NOR2_X1 i_0_643 (.ZN (\pp[13] [29] ), .A1 (n_0_50), .A2 (n_0_18));
NOR2_X1 i_0_642 (.ZN (\pp[13] [28] ), .A1 (n_0_50), .A2 (n_0_17));
NOR2_X1 i_0_641 (.ZN (\pp[13] [27] ), .A1 (n_0_50), .A2 (n_0_16));
NOR2_X1 i_0_640 (.ZN (\pp[13] [26] ), .A1 (n_0_50), .A2 (sgo__n50));
NOR2_X1 i_0_639 (.ZN (\pp[13] [25] ), .A1 (n_0_50), .A2 (sgo__n240));
NOR2_X1 i_0_638 (.ZN (\pp[13] [24] ), .A1 (n_0_50), .A2 (n_0_13));
NOR2_X1 i_0_637 (.ZN (\pp[13] [23] ), .A1 (n_0_50), .A2 (sgo__n157));
NOR2_X1 i_0_636 (.ZN (\pp[13] [22] ), .A1 (n_0_50), .A2 (sgo__n177));
NOR2_X1 i_0_635 (.ZN (\pp[13] [21] ), .A1 (n_0_50), .A2 (sgo__n162));
NOR2_X1 i_0_634 (.ZN (\pp[13] [20] ), .A1 (n_0_50), .A2 (n_0_9));
NOR2_X1 i_0_633 (.ZN (\pp[13] [19] ), .A1 (n_0_50), .A2 (sgo__n184));
NOR2_X1 i_0_632 (.ZN (\pp[13] [18] ), .A1 (n_0_50), .A2 (sgo__n172));
NOR2_X1 i_0_631 (.ZN (\pp[13] [17] ), .A1 (n_0_50), .A2 (sgo__n205));
NOR2_X1 i_0_630 (.ZN (\pp[13] [16] ), .A1 (n_0_50), .A2 (n_0_5));
NOR2_X1 i_0_629 (.ZN (\pp[13] [15] ), .A1 (n_0_50), .A2 (sgo__n66));
NOR2_X2 i_0_628 (.ZN (\pp[13] [14] ), .A1 (n_0_50), .A2 (sgo__n31));
NOR2_X1 i_0_627 (.ZN (\pp[13] [13] ), .A1 (n_0_50), .A2 (sgo__n39));
INV_X4 i_0_626 (.ZN (n_0_50), .A (x[13]));
NOR2_X1 i_0_625 (.ZN (\pp[14] [62] ), .A1 (n_0_49), .A2 (n_0_33));
NOR2_X1 i_0_624 (.ZN (\pp[14] [44] ), .A1 (n_0_49), .A2 (n_0_32));
NOR2_X1 i_0_623 (.ZN (\pp[14] [43] ), .A1 (n_0_49), .A2 (n_0_31));
NOR2_X1 i_0_622 (.ZN (\pp[14] [42] ), .A1 (n_0_49), .A2 (n_0_30));
NOR2_X1 i_0_621 (.ZN (\pp[14] [41] ), .A1 (n_0_49), .A2 (n_0_29));
NOR2_X1 i_0_620 (.ZN (\pp[14] [40] ), .A1 (n_0_49), .A2 (n_0_28));
NOR2_X1 i_0_619 (.ZN (\pp[14] [39] ), .A1 (n_0_49), .A2 (n_0_27));
NOR2_X1 i_0_618 (.ZN (\pp[14] [38] ), .A1 (n_0_49), .A2 (n_0_26));
NOR2_X1 i_0_617 (.ZN (\pp[14] [37] ), .A1 (n_0_49), .A2 (n_0_25));
NOR2_X1 i_0_616 (.ZN (\pp[14] [36] ), .A1 (n_0_49), .A2 (n_0_24));
NOR2_X1 i_0_615 (.ZN (\pp[14] [35] ), .A1 (n_0_49), .A2 (n_0_23));
NOR2_X1 i_0_614 (.ZN (\pp[14] [34] ), .A1 (n_0_49), .A2 (n_0_22));
NOR2_X1 i_0_613 (.ZN (\pp[14] [33] ), .A1 (n_0_49), .A2 (n_0_21));
NOR2_X1 i_0_612 (.ZN (\pp[14] [32] ), .A1 (n_0_49), .A2 (n_0_20));
NOR2_X1 i_0_611 (.ZN (\pp[14] [31] ), .A1 (n_0_49), .A2 (n_0_19));
NOR2_X1 i_0_610 (.ZN (\pp[14] [30] ), .A1 (n_0_49), .A2 (n_0_18));
NOR2_X1 i_0_609 (.ZN (\pp[14] [29] ), .A1 (n_0_49), .A2 (n_0_17));
NOR2_X1 i_0_608 (.ZN (\pp[14] [28] ), .A1 (n_0_49), .A2 (n_0_16));
NOR2_X1 i_0_607 (.ZN (\pp[14] [27] ), .A1 (n_0_49), .A2 (sgo__n50));
NOR2_X1 i_0_606 (.ZN (\pp[14] [26] ), .A1 (n_0_49), .A2 (sgo__n240));
NOR2_X1 i_0_605 (.ZN (\pp[14] [25] ), .A1 (n_0_49), .A2 (sgo__n106));
NOR2_X1 i_0_604 (.ZN (\pp[14] [24] ), .A1 (n_0_49), .A2 (sgo__n157));
NOR2_X1 i_0_603 (.ZN (\pp[14] [23] ), .A1 (n_0_49), .A2 (n_0_11));
NOR2_X1 i_0_602 (.ZN (\pp[14] [22] ), .A1 (n_0_49), .A2 (sgo__n162));
NOR2_X1 i_0_601 (.ZN (\pp[14] [21] ), .A1 (n_0_49), .A2 (n_0_9));
NOR2_X1 i_0_600 (.ZN (\pp[14] [20] ), .A1 (n_0_49), .A2 (sgo__n184));
NOR2_X1 i_0_599 (.ZN (\pp[14] [19] ), .A1 (n_0_49), .A2 (sgo__n172));
NOR2_X1 i_0_598 (.ZN (\pp[14] [18] ), .A1 (n_0_49), .A2 (sgo__n205));
NOR2_X1 i_0_597 (.ZN (\pp[14] [17] ), .A1 (n_0_49), .A2 (n_0_5));
NOR2_X2 i_0_596 (.ZN (\pp[14] [16] ), .A1 (n_0_49), .A2 (sgo__n66));
NOR2_X1 i_0_595 (.ZN (\pp[14] [15] ), .A1 (n_0_49), .A2 (sgo__n31));
NOR2_X2 i_0_594 (.ZN (\pp[14] [14] ), .A1 (n_0_49), .A2 (sgo__n39));
INV_X8 i_0_593 (.ZN (n_0_49), .A (x[14]));
NOR2_X1 i_0_592 (.ZN (\pp[15] [62] ), .A1 (n_0_48), .A2 (n_0_33));
NOR2_X1 i_0_591 (.ZN (\pp[15] [45] ), .A1 (n_0_48), .A2 (n_0_32));
NOR2_X1 i_0_590 (.ZN (\pp[15] [44] ), .A1 (n_0_48), .A2 (n_0_31));
NOR2_X1 i_0_589 (.ZN (\pp[15] [43] ), .A1 (n_0_48), .A2 (n_0_30));
NOR2_X1 i_0_588 (.ZN (\pp[15] [42] ), .A1 (n_0_48), .A2 (n_0_29));
NOR2_X1 i_0_587 (.ZN (\pp[15] [41] ), .A1 (n_0_48), .A2 (n_0_28));
NOR2_X1 i_0_586 (.ZN (\pp[15] [40] ), .A1 (n_0_48), .A2 (n_0_27));
NOR2_X1 i_0_585 (.ZN (\pp[15] [39] ), .A1 (n_0_48), .A2 (n_0_26));
NOR2_X1 i_0_584 (.ZN (\pp[15] [38] ), .A1 (n_0_48), .A2 (n_0_25));
NOR2_X1 i_0_583 (.ZN (\pp[15] [37] ), .A1 (n_0_48), .A2 (n_0_24));
NOR2_X1 i_0_582 (.ZN (\pp[15] [36] ), .A1 (n_0_48), .A2 (n_0_23));
NOR2_X1 i_0_581 (.ZN (\pp[15] [35] ), .A1 (n_0_48), .A2 (n_0_22));
NOR2_X1 i_0_580 (.ZN (\pp[15] [34] ), .A1 (n_0_48), .A2 (n_0_21));
NOR2_X1 i_0_579 (.ZN (\pp[15] [33] ), .A1 (n_0_48), .A2 (n_0_20));
NOR2_X1 i_0_578 (.ZN (\pp[15] [32] ), .A1 (n_0_48), .A2 (n_0_19));
NOR2_X1 i_0_577 (.ZN (\pp[15] [31] ), .A1 (n_0_48), .A2 (n_0_18));
NOR2_X1 i_0_576 (.ZN (\pp[15] [30] ), .A1 (n_0_48), .A2 (n_0_17));
NOR2_X1 i_0_575 (.ZN (\pp[15] [29] ), .A1 (n_0_48), .A2 (n_0_16));
NOR2_X1 i_0_574 (.ZN (\pp[15] [28] ), .A1 (n_0_48), .A2 (sgo__n50));
NOR2_X1 i_0_573 (.ZN (\pp[15] [27] ), .A1 (n_0_48), .A2 (sgo__n240));
NOR2_X1 i_0_572 (.ZN (\pp[15] [26] ), .A1 (n_0_48), .A2 (sgo__n106));
NOR2_X1 i_0_571 (.ZN (\pp[15] [25] ), .A1 (n_0_48), .A2 (sgo__n157));
NOR2_X1 i_0_570 (.ZN (\pp[15] [24] ), .A1 (n_0_48), .A2 (sgo__n177));
NOR2_X1 i_0_569 (.ZN (\pp[15] [23] ), .A1 (n_0_48), .A2 (sgo__n162));
NOR2_X1 i_0_568 (.ZN (\pp[15] [22] ), .A1 (n_0_48), .A2 (sgo__n74));
NOR2_X1 i_0_567 (.ZN (\pp[15] [21] ), .A1 (n_0_48), .A2 (sgo__n184));
NOR2_X1 i_0_566 (.ZN (\pp[15] [20] ), .A1 (n_0_48), .A2 (sgo__n172));
NOR2_X1 i_0_565 (.ZN (\pp[15] [19] ), .A1 (n_0_48), .A2 (sgo__n205));
NOR2_X1 i_0_564 (.ZN (\pp[15] [18] ), .A1 (n_0_48), .A2 (n_0_5));
NOR2_X1 i_0_563 (.ZN (\pp[15] [17] ), .A1 (n_0_48), .A2 (sgo__n69));
NOR2_X1 i_0_562 (.ZN (\pp[15] [16] ), .A1 (n_0_48), .A2 (sgo__n31));
NOR2_X1 i_0_561 (.ZN (\pp[15] [15] ), .A1 (n_0_48), .A2 (sgo__n39));
INV_X4 i_0_560 (.ZN (n_0_48), .A (x[15]));
NOR2_X1 i_0_559 (.ZN (\pp[16] [62] ), .A1 (n_0_47), .A2 (n_0_33));
NOR2_X1 i_0_558 (.ZN (\pp[16] [46] ), .A1 (n_0_47), .A2 (n_0_32));
NOR2_X1 i_0_557 (.ZN (\pp[16] [45] ), .A1 (n_0_47), .A2 (n_0_31));
NOR2_X1 i_0_556 (.ZN (\pp[16] [44] ), .A1 (n_0_47), .A2 (n_0_30));
NOR2_X1 i_0_555 (.ZN (\pp[16] [43] ), .A1 (n_0_47), .A2 (n_0_29));
NOR2_X1 i_0_554 (.ZN (\pp[16] [42] ), .A1 (n_0_47), .A2 (n_0_28));
NOR2_X1 i_0_553 (.ZN (\pp[16] [41] ), .A1 (n_0_47), .A2 (n_0_27));
NOR2_X1 i_0_552 (.ZN (\pp[16] [40] ), .A1 (n_0_47), .A2 (n_0_26));
NOR2_X1 i_0_551 (.ZN (\pp[16] [39] ), .A1 (n_0_47), .A2 (n_0_25));
NOR2_X1 i_0_550 (.ZN (\pp[16] [38] ), .A1 (n_0_47), .A2 (n_0_24));
NOR2_X1 i_0_549 (.ZN (\pp[16] [37] ), .A1 (n_0_47), .A2 (n_0_23));
NOR2_X1 i_0_548 (.ZN (\pp[16] [36] ), .A1 (n_0_47), .A2 (n_0_22));
NOR2_X1 i_0_547 (.ZN (\pp[16] [35] ), .A1 (n_0_47), .A2 (n_0_21));
NOR2_X1 i_0_546 (.ZN (\pp[16] [34] ), .A1 (n_0_47), .A2 (n_0_20));
NOR2_X1 i_0_545 (.ZN (\pp[16] [33] ), .A1 (n_0_47), .A2 (n_0_19));
NOR2_X1 i_0_544 (.ZN (\pp[16] [32] ), .A1 (n_0_47), .A2 (n_0_18));
NOR2_X1 i_0_543 (.ZN (\pp[16] [31] ), .A1 (n_0_47), .A2 (n_0_17));
NOR2_X1 i_0_542 (.ZN (\pp[16] [30] ), .A1 (n_0_47), .A2 (n_0_16));
NOR2_X1 i_0_541 (.ZN (\pp[16] [29] ), .A1 (n_0_47), .A2 (sgo__n50));
NOR2_X1 i_0_540 (.ZN (\pp[16] [28] ), .A1 (n_0_47), .A2 (sgo__n240));
NOR2_X1 i_0_539 (.ZN (\pp[16] [27] ), .A1 (n_0_47), .A2 (sgo__n106));
NOR2_X1 i_0_538 (.ZN (\pp[16] [26] ), .A1 (n_0_47), .A2 (sgo__n157));
NOR2_X1 i_0_537 (.ZN (\pp[16] [25] ), .A1 (n_0_47), .A2 (sgo__n133));
NOR2_X1 i_0_536 (.ZN (\pp[16] [24] ), .A1 (n_0_47), .A2 (sgo__n162));
NOR2_X1 i_0_535 (.ZN (\pp[16] [23] ), .A1 (n_0_47), .A2 (sgo__n74));
NOR2_X1 i_0_534 (.ZN (\pp[16] [22] ), .A1 (n_0_47), .A2 (sgo__n184));
NOR2_X1 i_0_533 (.ZN (\pp[16] [21] ), .A1 (n_0_47), .A2 (sgo__n172));
NOR2_X1 i_0_532 (.ZN (\pp[16] [20] ), .A1 (n_0_47), .A2 (sgo__n205));
NOR2_X1 i_0_531 (.ZN (\pp[16] [19] ), .A1 (n_0_47), .A2 (n_0_5));
NOR2_X1 i_0_530 (.ZN (\pp[16] [18] ), .A1 (n_0_47), .A2 (sgo__n69));
NOR2_X1 i_0_529 (.ZN (\pp[16] [17] ), .A1 (n_0_47), .A2 (sgo__n31));
NOR2_X1 i_0_528 (.ZN (\pp[16] [16] ), .A1 (n_0_47), .A2 (sgo__n39));
INV_X4 i_0_527 (.ZN (n_0_47), .A (x[16]));
NOR2_X1 i_0_526 (.ZN (\pp[17] [62] ), .A1 (n_0_46), .A2 (n_0_33));
NOR2_X1 i_0_525 (.ZN (\pp[17] [47] ), .A1 (n_0_46), .A2 (n_0_32));
NOR2_X1 i_0_524 (.ZN (\pp[17] [46] ), .A1 (n_0_46), .A2 (n_0_31));
NOR2_X1 i_0_523 (.ZN (\pp[17] [45] ), .A1 (n_0_46), .A2 (n_0_30));
NOR2_X1 i_0_522 (.ZN (\pp[17] [44] ), .A1 (n_0_46), .A2 (n_0_29));
NOR2_X1 i_0_521 (.ZN (\pp[17] [43] ), .A1 (n_0_46), .A2 (n_0_28));
NOR2_X1 i_0_520 (.ZN (\pp[17] [42] ), .A1 (n_0_46), .A2 (n_0_27));
NOR2_X1 i_0_519 (.ZN (\pp[17] [41] ), .A1 (n_0_46), .A2 (n_0_26));
NOR2_X1 i_0_518 (.ZN (\pp[17] [40] ), .A1 (n_0_46), .A2 (n_0_25));
NOR2_X1 i_0_517 (.ZN (\pp[17] [39] ), .A1 (n_0_46), .A2 (n_0_24));
NOR2_X1 i_0_516 (.ZN (\pp[17] [38] ), .A1 (n_0_46), .A2 (n_0_23));
NOR2_X1 i_0_515 (.ZN (\pp[17] [37] ), .A1 (n_0_46), .A2 (n_0_22));
NOR2_X1 i_0_514 (.ZN (\pp[17] [36] ), .A1 (n_0_46), .A2 (n_0_21));
NOR2_X1 i_0_513 (.ZN (\pp[17] [35] ), .A1 (n_0_46), .A2 (n_0_20));
NOR2_X1 i_0_512 (.ZN (\pp[17] [34] ), .A1 (n_0_46), .A2 (n_0_19));
NOR2_X1 i_0_511 (.ZN (\pp[17] [33] ), .A1 (n_0_46), .A2 (n_0_18));
NOR2_X1 i_0_510 (.ZN (\pp[17] [32] ), .A1 (n_0_46), .A2 (n_0_17));
NOR2_X1 i_0_509 (.ZN (\pp[17] [31] ), .A1 (n_0_46), .A2 (n_0_16));
NOR2_X1 i_0_508 (.ZN (\pp[17] [30] ), .A1 (n_0_46), .A2 (sgo__n50));
NOR2_X1 i_0_507 (.ZN (\pp[17] [29] ), .A1 (n_0_46), .A2 (sgo__n140));
NOR2_X1 i_0_506 (.ZN (\pp[17] [28] ), .A1 (n_0_46), .A2 (sgo__n106));
NOR2_X1 i_0_505 (.ZN (\pp[17] [27] ), .A1 (n_0_46), .A2 (sgo__n157));
NOR2_X1 i_0_504 (.ZN (\pp[17] [26] ), .A1 (n_0_46), .A2 (sgo__n133));
NOR2_X1 i_0_503 (.ZN (\pp[17] [25] ), .A1 (n_0_46), .A2 (sgo__n162));
NOR2_X1 i_0_502 (.ZN (\pp[17] [24] ), .A1 (n_0_46), .A2 (sgo__n74));
NOR2_X1 i_0_501 (.ZN (\pp[17] [23] ), .A1 (n_0_46), .A2 (sgo__n184));
NOR2_X1 i_0_500 (.ZN (\pp[17] [22] ), .A1 (n_0_46), .A2 (sgo__n172));
NOR2_X1 i_0_499 (.ZN (\pp[17] [21] ), .A1 (n_0_46), .A2 (sgo__n205));
NOR2_X1 i_0_498 (.ZN (\pp[17] [20] ), .A1 (n_0_46), .A2 (n_0_5));
NOR2_X1 i_0_497 (.ZN (\pp[17] [19] ), .A1 (n_0_46), .A2 (sgo__n69));
NOR2_X1 i_0_496 (.ZN (\pp[17] [18] ), .A1 (n_0_46), .A2 (sgo__n31));
NOR2_X1 i_0_495 (.ZN (\pp[17] [17] ), .A1 (n_0_46), .A2 (sgo__n39));
INV_X4 i_0_494 (.ZN (n_0_46), .A (x[17]));
NOR2_X1 i_0_493 (.ZN (\pp[18] [63] ), .A1 (n_0_45), .A2 (n_0_33));
NOR2_X1 i_0_492 (.ZN (\pp[18] [48] ), .A1 (n_0_45), .A2 (n_0_32));
NOR2_X1 i_0_491 (.ZN (\pp[18] [47] ), .A1 (n_0_45), .A2 (n_0_31));
NOR2_X1 i_0_490 (.ZN (\pp[18] [46] ), .A1 (n_0_45), .A2 (n_0_30));
NOR2_X1 i_0_489 (.ZN (\pp[18] [45] ), .A1 (n_0_45), .A2 (n_0_29));
NOR2_X1 i_0_488 (.ZN (\pp[18] [44] ), .A1 (n_0_45), .A2 (n_0_28));
NOR2_X1 i_0_487 (.ZN (\pp[18] [43] ), .A1 (n_0_45), .A2 (n_0_27));
NOR2_X1 i_0_486 (.ZN (\pp[18] [42] ), .A1 (n_0_45), .A2 (n_0_26));
NOR2_X1 i_0_485 (.ZN (\pp[18] [41] ), .A1 (n_0_45), .A2 (n_0_25));
NOR2_X1 i_0_484 (.ZN (\pp[18] [40] ), .A1 (n_0_45), .A2 (n_0_24));
NOR2_X1 i_0_483 (.ZN (\pp[18] [39] ), .A1 (n_0_45), .A2 (n_0_23));
NOR2_X1 i_0_482 (.ZN (\pp[18] [38] ), .A1 (n_0_45), .A2 (n_0_22));
NOR2_X1 i_0_481 (.ZN (\pp[18] [37] ), .A1 (n_0_45), .A2 (n_0_21));
NOR2_X1 i_0_480 (.ZN (\pp[18] [36] ), .A1 (n_0_45), .A2 (n_0_20));
NOR2_X1 i_0_479 (.ZN (\pp[18] [35] ), .A1 (n_0_45), .A2 (n_0_19));
NOR2_X1 i_0_478 (.ZN (\pp[18] [34] ), .A1 (n_0_45), .A2 (n_0_18));
NOR2_X1 i_0_477 (.ZN (\pp[18] [33] ), .A1 (n_0_45), .A2 (n_0_17));
NOR2_X1 i_0_476 (.ZN (\pp[18] [32] ), .A1 (n_0_45), .A2 (n_0_16));
NOR2_X1 i_0_475 (.ZN (\pp[18] [31] ), .A1 (n_0_45), .A2 (sgo__n50));
NOR2_X1 i_0_474 (.ZN (\pp[18] [30] ), .A1 (n_0_45), .A2 (sgo__n140));
NOR2_X1 i_0_473 (.ZN (\pp[18] [29] ), .A1 (n_0_45), .A2 (sgo__n106));
NOR2_X1 i_0_472 (.ZN (\pp[18] [28] ), .A1 (n_0_45), .A2 (sgo__n157));
NOR2_X1 i_0_471 (.ZN (\pp[18] [27] ), .A1 (n_0_45), .A2 (sgo__n133));
NOR2_X1 i_0_470 (.ZN (\pp[18] [26] ), .A1 (n_0_45), .A2 (sgo__n162));
NOR2_X1 i_0_469 (.ZN (\pp[18] [25] ), .A1 (n_0_45), .A2 (sgo__n74));
NOR2_X1 i_0_468 (.ZN (\pp[18] [24] ), .A1 (n_0_45), .A2 (sgo__n184));
NOR2_X1 i_0_467 (.ZN (\pp[18] [23] ), .A1 (n_0_45), .A2 (sgo__n172));
NOR2_X1 i_0_466 (.ZN (\pp[18] [22] ), .A1 (n_0_45), .A2 (sgo__n205));
NOR2_X1 i_0_465 (.ZN (\pp[18] [21] ), .A1 (n_0_45), .A2 (n_0_5));
NOR2_X1 i_0_464 (.ZN (\pp[18] [20] ), .A1 (n_0_45), .A2 (sgo__n69));
NOR2_X1 i_0_463 (.ZN (\pp[18] [19] ), .A1 (n_0_45), .A2 (sgo__n31));
NOR2_X1 i_0_462 (.ZN (\pp[18] [18] ), .A1 (n_0_45), .A2 (sgo__n39));
INV_X4 i_0_461 (.ZN (n_0_45), .A (x[18]));
NOR2_X1 i_0_460 (.ZN (\pp[19] [63] ), .A1 (n_0_44), .A2 (n_0_33));
NOR2_X1 i_0_459 (.ZN (\pp[19] [49] ), .A1 (n_0_44), .A2 (n_0_32));
NOR2_X1 i_0_458 (.ZN (\pp[19] [48] ), .A1 (n_0_44), .A2 (n_0_31));
NOR2_X1 i_0_457 (.ZN (\pp[19] [47] ), .A1 (n_0_44), .A2 (n_0_30));
NOR2_X1 i_0_456 (.ZN (\pp[19] [46] ), .A1 (n_0_44), .A2 (n_0_29));
NOR2_X1 i_0_455 (.ZN (\pp[19] [45] ), .A1 (n_0_44), .A2 (n_0_28));
NOR2_X1 i_0_454 (.ZN (\pp[19] [44] ), .A1 (n_0_44), .A2 (n_0_27));
NOR2_X1 i_0_453 (.ZN (\pp[19] [43] ), .A1 (n_0_44), .A2 (n_0_26));
NOR2_X1 i_0_452 (.ZN (\pp[19] [42] ), .A1 (n_0_44), .A2 (n_0_25));
NOR2_X1 i_0_451 (.ZN (\pp[19] [41] ), .A1 (n_0_44), .A2 (n_0_24));
NOR2_X1 i_0_450 (.ZN (\pp[19] [40] ), .A1 (n_0_44), .A2 (n_0_23));
NOR2_X1 i_0_449 (.ZN (\pp[19] [39] ), .A1 (n_0_44), .A2 (n_0_22));
NOR2_X1 i_0_448 (.ZN (\pp[19] [38] ), .A1 (n_0_44), .A2 (n_0_21));
NOR2_X1 i_0_447 (.ZN (\pp[19] [37] ), .A1 (n_0_44), .A2 (n_0_20));
NOR2_X1 i_0_446 (.ZN (\pp[19] [36] ), .A1 (n_0_44), .A2 (n_0_19));
NOR2_X1 i_0_445 (.ZN (\pp[19] [35] ), .A1 (n_0_44), .A2 (n_0_18));
NOR2_X1 i_0_444 (.ZN (\pp[19] [34] ), .A1 (n_0_44), .A2 (n_0_17));
NOR2_X1 i_0_443 (.ZN (\pp[19] [33] ), .A1 (n_0_44), .A2 (n_0_16));
NOR2_X1 i_0_442 (.ZN (\pp[19] [32] ), .A1 (n_0_44), .A2 (sgo__n50));
NOR2_X1 i_0_441 (.ZN (\pp[19] [31] ), .A1 (n_0_44), .A2 (sgo__n240));
NOR2_X1 i_0_440 (.ZN (\pp[19] [30] ), .A1 (n_0_44), .A2 (sgo__n106));
NOR2_X1 i_0_439 (.ZN (\pp[19] [29] ), .A1 (n_0_44), .A2 (sgo__n157));
NOR2_X1 i_0_438 (.ZN (\pp[19] [28] ), .A1 (n_0_44), .A2 (sgo__n133));
NOR2_X1 i_0_437 (.ZN (\pp[19] [27] ), .A1 (n_0_44), .A2 (sgo__n162));
NOR2_X1 i_0_436 (.ZN (\pp[19] [26] ), .A1 (n_0_44), .A2 (sgo__n74));
NOR2_X1 i_0_435 (.ZN (\pp[19] [25] ), .A1 (n_0_44), .A2 (sgo__n184));
NOR2_X1 i_0_434 (.ZN (\pp[19] [24] ), .A1 (n_0_44), .A2 (sgo__n172));
NOR2_X1 i_0_433 (.ZN (\pp[19] [23] ), .A1 (n_0_44), .A2 (n_0_6));
NOR2_X1 i_0_432 (.ZN (\pp[19] [22] ), .A1 (n_0_44), .A2 (n_0_5));
NOR2_X1 i_0_431 (.ZN (\pp[19] [21] ), .A1 (n_0_44), .A2 (sgo__n69));
NOR2_X1 i_0_430 (.ZN (\pp[19] [20] ), .A1 (n_0_44), .A2 (sgo__n31));
NOR2_X1 i_0_429 (.ZN (\pp[19] [19] ), .A1 (n_0_44), .A2 (sgo__n39));
INV_X4 i_0_428 (.ZN (n_0_44), .A (x[19]));
NOR2_X1 i_0_427 (.ZN (\pp[20] [63] ), .A1 (n_0_43), .A2 (n_0_33));
NOR2_X1 i_0_426 (.ZN (\pp[20] [50] ), .A1 (n_0_43), .A2 (n_0_32));
NOR2_X1 i_0_425 (.ZN (\pp[20] [49] ), .A1 (n_0_43), .A2 (n_0_31));
NOR2_X1 i_0_424 (.ZN (\pp[20] [48] ), .A1 (n_0_43), .A2 (n_0_30));
NOR2_X1 i_0_423 (.ZN (\pp[20] [47] ), .A1 (n_0_43), .A2 (n_0_29));
NOR2_X1 i_0_422 (.ZN (\pp[20] [46] ), .A1 (drc_ipo_n910), .A2 (n_0_28));
NOR2_X1 i_0_421 (.ZN (\pp[20] [45] ), .A1 (drc_ipo_n910), .A2 (n_0_27));
NOR2_X1 i_0_420 (.ZN (\pp[20] [44] ), .A1 (drc_ipo_n910), .A2 (n_0_26));
NOR2_X1 i_0_419 (.ZN (\pp[20] [43] ), .A1 (drc_ipo_n910), .A2 (n_0_25));
NOR2_X1 i_0_418 (.ZN (\pp[20] [42] ), .A1 (drc_ipo_n910), .A2 (n_0_24));
NOR2_X1 i_0_417 (.ZN (\pp[20] [41] ), .A1 (drc_ipo_n910), .A2 (n_0_23));
NOR2_X1 i_0_416 (.ZN (\pp[20] [40] ), .A1 (drc_ipo_n910), .A2 (n_0_22));
NOR2_X1 i_0_415 (.ZN (\pp[20] [39] ), .A1 (drc_ipo_n910), .A2 (n_0_21));
NOR2_X1 i_0_414 (.ZN (\pp[20] [38] ), .A1 (drc_ipo_n910), .A2 (n_0_20));
NOR2_X1 i_0_413 (.ZN (\pp[20] [37] ), .A1 (drc_ipo_n910), .A2 (n_0_19));
NOR2_X1 i_0_412 (.ZN (\pp[20] [36] ), .A1 (drc_ipo_n910), .A2 (n_0_18));
NOR2_X1 i_0_411 (.ZN (\pp[20] [35] ), .A1 (drc_ipo_n910), .A2 (n_0_17));
NOR2_X1 i_0_410 (.ZN (\pp[20] [34] ), .A1 (drc_ipo_n910), .A2 (n_0_16));
NOR2_X1 i_0_409 (.ZN (\pp[20] [33] ), .A1 (drc_ipo_n910), .A2 (sgo__n50));
NOR2_X1 i_0_408 (.ZN (\pp[20] [32] ), .A1 (drc_ipo_n910), .A2 (sgo__n240));
NOR2_X1 i_0_407 (.ZN (\pp[20] [31] ), .A1 (drc_ipo_n910), .A2 (sgo__n106));
NOR2_X1 i_0_406 (.ZN (\pp[20] [30] ), .A1 (drc_ipo_n910), .A2 (sgo__n157));
NOR2_X1 i_0_405 (.ZN (\pp[20] [29] ), .A1 (drc_ipo_n910), .A2 (sgo__n133));
NOR2_X1 i_0_404 (.ZN (\pp[20] [28] ), .A1 (drc_ipo_n910), .A2 (sgo__n162));
NOR2_X1 i_0_403 (.ZN (\pp[20] [27] ), .A1 (drc_ipo_n910), .A2 (sgo__n74));
NOR2_X1 i_0_402 (.ZN (\pp[20] [26] ), .A1 (drc_ipo_n910), .A2 (sgo__n184));
NOR2_X1 i_0_401 (.ZN (\pp[20] [25] ), .A1 (drc_ipo_n910), .A2 (sgo__n172));
NOR2_X1 i_0_400 (.ZN (\pp[20] [24] ), .A1 (drc_ipo_n910), .A2 (n_0_6));
NOR2_X1 i_0_399 (.ZN (\pp[20] [23] ), .A1 (drc_ipo_n910), .A2 (n_0_5));
NOR2_X1 i_0_398 (.ZN (\pp[20] [22] ), .A1 (drc_ipo_n910), .A2 (n_0_4));
NOR2_X1 i_0_397 (.ZN (\pp[20] [21] ), .A1 (n_0_43), .A2 (sgo__n34));
NOR2_X1 i_0_396 (.ZN (\pp[20] [20] ), .A1 (n_0_43), .A2 (n_0_2));
INV_X4 i_0_395 (.ZN (n_0_43), .A (x[20]));
NOR2_X1 i_0_394 (.ZN (\pp[21] [63] ), .A1 (n_0_42), .A2 (n_0_33));
NOR2_X1 i_0_393 (.ZN (\pp[21] [51] ), .A1 (n_0_42), .A2 (n_0_32));
NOR2_X1 i_0_392 (.ZN (\pp[21] [50] ), .A1 (n_0_42), .A2 (n_0_31));
NOR2_X1 i_0_391 (.ZN (\pp[21] [49] ), .A1 (n_0_42), .A2 (n_0_30));
NOR2_X1 i_0_390 (.ZN (\pp[21] [48] ), .A1 (drc_ipo_n911), .A2 (n_0_29));
NOR2_X1 i_0_389 (.ZN (\pp[21] [47] ), .A1 (drc_ipo_n911), .A2 (n_0_28));
NOR2_X1 i_0_388 (.ZN (\pp[21] [46] ), .A1 (drc_ipo_n911), .A2 (n_0_27));
NOR2_X1 i_0_387 (.ZN (\pp[21] [45] ), .A1 (drc_ipo_n911), .A2 (n_0_26));
NOR2_X1 i_0_386 (.ZN (\pp[21] [44] ), .A1 (drc_ipo_n911), .A2 (n_0_25));
NOR2_X1 i_0_385 (.ZN (\pp[21] [43] ), .A1 (drc_ipo_n911), .A2 (n_0_24));
NOR2_X1 i_0_384 (.ZN (\pp[21] [42] ), .A1 (drc_ipo_n911), .A2 (n_0_23));
NOR2_X1 i_0_383 (.ZN (\pp[21] [41] ), .A1 (drc_ipo_n911), .A2 (n_0_22));
NOR2_X1 i_0_382 (.ZN (\pp[21] [40] ), .A1 (drc_ipo_n911), .A2 (n_0_21));
NOR2_X1 i_0_381 (.ZN (\pp[21] [39] ), .A1 (drc_ipo_n911), .A2 (n_0_20));
NOR2_X1 i_0_380 (.ZN (\pp[21] [38] ), .A1 (drc_ipo_n911), .A2 (n_0_19));
NOR2_X1 i_0_379 (.ZN (\pp[21] [37] ), .A1 (drc_ipo_n911), .A2 (n_0_18));
NOR2_X1 i_0_378 (.ZN (\pp[21] [36] ), .A1 (drc_ipo_n911), .A2 (n_0_17));
NOR2_X1 i_0_377 (.ZN (\pp[21] [35] ), .A1 (drc_ipo_n911), .A2 (n_0_16));
NOR2_X1 i_0_376 (.ZN (\pp[21] [34] ), .A1 (drc_ipo_n911), .A2 (sgo__n50));
NOR2_X1 i_0_375 (.ZN (\pp[21] [33] ), .A1 (drc_ipo_n911), .A2 (sgo__n240));
NOR2_X1 i_0_374 (.ZN (\pp[21] [32] ), .A1 (drc_ipo_n911), .A2 (sgo__n106));
NOR2_X1 i_0_373 (.ZN (\pp[21] [31] ), .A1 (drc_ipo_n911), .A2 (sgo__n157));
NOR2_X1 i_0_372 (.ZN (\pp[21] [30] ), .A1 (drc_ipo_n911), .A2 (sgo__n133));
NOR2_X1 i_0_371 (.ZN (\pp[21] [29] ), .A1 (drc_ipo_n911), .A2 (sgo__n162));
NOR2_X1 i_0_370 (.ZN (\pp[21] [28] ), .A1 (drc_ipo_n911), .A2 (sgo__n74));
NOR2_X1 i_0_369 (.ZN (\pp[21] [27] ), .A1 (drc_ipo_n911), .A2 (sgo__n184));
NOR2_X1 i_0_368 (.ZN (\pp[21] [26] ), .A1 (drc_ipo_n911), .A2 (sgo__n172));
NOR2_X1 i_0_367 (.ZN (\pp[21] [25] ), .A1 (drc_ipo_n911), .A2 (n_0_6));
NOR2_X1 i_0_366 (.ZN (\pp[21] [24] ), .A1 (drc_ipo_n911), .A2 (n_0_5));
NOR2_X1 i_0_365 (.ZN (\pp[21] [23] ), .A1 (drc_ipo_n911), .A2 (n_0_4));
NOR2_X1 i_0_364 (.ZN (\pp[21] [22] ), .A1 (n_0_42), .A2 (sgo__n34));
NOR2_X1 i_0_363 (.ZN (\pp[21] [21] ), .A1 (n_0_42), .A2 (n_0_2));
INV_X4 i_0_362 (.ZN (n_0_42), .A (x[21]));
NOR2_X1 i_0_361 (.ZN (\pp[22] [63] ), .A1 (n_0_41), .A2 (n_0_33));
NOR2_X1 i_0_360 (.ZN (\pp[22] [52] ), .A1 (n_0_41), .A2 (n_0_32));
NOR2_X1 i_0_359 (.ZN (\pp[22] [51] ), .A1 (n_0_41), .A2 (n_0_31));
NOR2_X1 i_0_358 (.ZN (\pp[22] [50] ), .A1 (n_0_41), .A2 (n_0_30));
NOR2_X1 i_0_357 (.ZN (\pp[22] [49] ), .A1 (n_0_41), .A2 (n_0_29));
NOR2_X1 i_0_356 (.ZN (\pp[22] [48] ), .A1 (n_0_41), .A2 (n_0_28));
NOR2_X1 i_0_355 (.ZN (\pp[22] [47] ), .A1 (n_0_41), .A2 (n_0_27));
NOR2_X1 i_0_354 (.ZN (\pp[22] [46] ), .A1 (n_0_41), .A2 (n_0_26));
NOR2_X1 i_0_353 (.ZN (\pp[22] [45] ), .A1 (n_0_41), .A2 (n_0_25));
NOR2_X1 i_0_352 (.ZN (\pp[22] [44] ), .A1 (n_0_41), .A2 (n_0_24));
NOR2_X1 i_0_351 (.ZN (\pp[22] [43] ), .A1 (n_0_41), .A2 (n_0_23));
NOR2_X1 i_0_350 (.ZN (\pp[22] [42] ), .A1 (n_0_41), .A2 (n_0_22));
NOR2_X1 i_0_349 (.ZN (\pp[22] [41] ), .A1 (n_0_41), .A2 (n_0_21));
NOR2_X1 i_0_348 (.ZN (\pp[22] [40] ), .A1 (n_0_41), .A2 (n_0_20));
NOR2_X1 i_0_347 (.ZN (\pp[22] [39] ), .A1 (n_0_41), .A2 (n_0_19));
NOR2_X1 i_0_346 (.ZN (\pp[22] [38] ), .A1 (n_0_41), .A2 (n_0_18));
NOR2_X1 i_0_345 (.ZN (\pp[22] [37] ), .A1 (n_0_41), .A2 (n_0_17));
NOR2_X1 i_0_344 (.ZN (\pp[22] [36] ), .A1 (n_0_41), .A2 (n_0_16));
NOR2_X1 i_0_343 (.ZN (\pp[22] [35] ), .A1 (n_0_41), .A2 (sgo__n50));
NOR2_X1 i_0_342 (.ZN (\pp[22] [34] ), .A1 (n_0_41), .A2 (sgo__n240));
NOR2_X1 i_0_341 (.ZN (\pp[22] [33] ), .A1 (n_0_41), .A2 (sgo__n106));
NOR2_X1 i_0_340 (.ZN (\pp[22] [32] ), .A1 (n_0_41), .A2 (sgo__n157));
NOR2_X1 i_0_339 (.ZN (\pp[22] [31] ), .A1 (n_0_41), .A2 (sgo__n133));
NOR2_X1 i_0_338 (.ZN (\pp[22] [30] ), .A1 (n_0_41), .A2 (sgo__n162));
NOR2_X1 i_0_337 (.ZN (\pp[22] [29] ), .A1 (n_0_41), .A2 (sgo__n74));
NOR2_X1 i_0_336 (.ZN (\pp[22] [28] ), .A1 (n_0_41), .A2 (sgo__n184));
NOR2_X1 i_0_335 (.ZN (\pp[22] [27] ), .A1 (n_0_41), .A2 (sgo__n172));
NOR2_X1 i_0_334 (.ZN (\pp[22] [26] ), .A1 (n_0_41), .A2 (sgo__n147));
NOR2_X1 i_0_333 (.ZN (\pp[22] [25] ), .A1 (n_0_41), .A2 (n_0_5));
NOR2_X1 i_0_332 (.ZN (\pp[22] [24] ), .A1 (n_0_41), .A2 (n_0_4));
NOR2_X1 i_0_331 (.ZN (\pp[22] [23] ), .A1 (n_0_41), .A2 (sgo__n34));
NOR2_X1 i_0_330 (.ZN (\pp[22] [22] ), .A1 (n_0_41), .A2 (n_0_2));
INV_X4 i_0_329 (.ZN (n_0_41), .A (x[22]));
NOR2_X1 i_0_328 (.ZN (\pp[23] [63] ), .A1 (n_0_40), .A2 (n_0_33));
NOR2_X1 i_0_327 (.ZN (\pp[23] [53] ), .A1 (n_0_40), .A2 (n_0_32));
NOR2_X1 i_0_326 (.ZN (\pp[23] [52] ), .A1 (n_0_40), .A2 (n_0_31));
NOR2_X1 i_0_325 (.ZN (\pp[23] [51] ), .A1 (n_0_40), .A2 (n_0_30));
NOR2_X1 i_0_324 (.ZN (\pp[23] [50] ), .A1 (n_0_40), .A2 (n_0_29));
NOR2_X1 i_0_323 (.ZN (\pp[23] [49] ), .A1 (n_0_40), .A2 (n_0_28));
NOR2_X1 i_0_322 (.ZN (\pp[23] [48] ), .A1 (n_0_40), .A2 (n_0_27));
NOR2_X1 i_0_321 (.ZN (\pp[23] [47] ), .A1 (n_0_40), .A2 (n_0_26));
NOR2_X1 i_0_320 (.ZN (\pp[23] [46] ), .A1 (n_0_40), .A2 (n_0_25));
NOR2_X1 i_0_319 (.ZN (\pp[23] [45] ), .A1 (n_0_40), .A2 (n_0_24));
NOR2_X1 i_0_318 (.ZN (\pp[23] [44] ), .A1 (n_0_40), .A2 (n_0_23));
NOR2_X1 i_0_317 (.ZN (\pp[23] [43] ), .A1 (n_0_40), .A2 (n_0_22));
NOR2_X1 i_0_316 (.ZN (\pp[23] [42] ), .A1 (n_0_40), .A2 (n_0_21));
NOR2_X1 i_0_315 (.ZN (\pp[23] [41] ), .A1 (n_0_40), .A2 (n_0_20));
NOR2_X1 i_0_314 (.ZN (\pp[23] [40] ), .A1 (n_0_40), .A2 (n_0_19));
NOR2_X1 i_0_313 (.ZN (\pp[23] [39] ), .A1 (n_0_40), .A2 (n_0_18));
NOR2_X1 i_0_312 (.ZN (\pp[23] [38] ), .A1 (n_0_40), .A2 (n_0_17));
NOR2_X1 i_0_311 (.ZN (\pp[23] [37] ), .A1 (n_0_40), .A2 (n_0_16));
NOR2_X1 i_0_310 (.ZN (\pp[23] [36] ), .A1 (n_0_40), .A2 (sgo__n50));
NOR2_X1 i_0_309 (.ZN (\pp[23] [35] ), .A1 (n_0_40), .A2 (sgo__n240));
NOR2_X1 i_0_308 (.ZN (\pp[23] [34] ), .A1 (n_0_40), .A2 (sgo__n106));
NOR2_X1 i_0_307 (.ZN (\pp[23] [33] ), .A1 (n_0_40), .A2 (sgo__n157));
NOR2_X1 i_0_306 (.ZN (\pp[23] [32] ), .A1 (n_0_40), .A2 (sgo__n133));
NOR2_X1 i_0_305 (.ZN (\pp[23] [31] ), .A1 (n_0_40), .A2 (sgo__n162));
NOR2_X1 i_0_304 (.ZN (\pp[23] [30] ), .A1 (n_0_40), .A2 (sgo__n74));
NOR2_X1 i_0_303 (.ZN (\pp[23] [29] ), .A1 (n_0_40), .A2 (sgo__n184));
NOR2_X1 i_0_302 (.ZN (\pp[23] [28] ), .A1 (n_0_40), .A2 (sgo__n172));
NOR2_X1 i_0_301 (.ZN (\pp[23] [27] ), .A1 (n_0_40), .A2 (sgo__n147));
NOR2_X1 i_0_300 (.ZN (\pp[23] [26] ), .A1 (n_0_40), .A2 (n_0_5));
NOR2_X1 i_0_299 (.ZN (\pp[23] [25] ), .A1 (n_0_40), .A2 (n_0_4));
NOR2_X1 i_0_298 (.ZN (\pp[23] [24] ), .A1 (n_0_40), .A2 (sgo__n34));
NOR2_X1 i_0_297 (.ZN (\pp[23] [23] ), .A1 (n_0_40), .A2 (n_0_2));
INV_X4 i_0_296 (.ZN (n_0_40), .A (x[23]));
NOR2_X1 i_0_295 (.ZN (\pp[24] [63] ), .A1 (n_0_39), .A2 (n_0_33));
NOR2_X1 i_0_294 (.ZN (\pp[24] [54] ), .A1 (n_0_39), .A2 (n_0_32));
NOR2_X1 i_0_293 (.ZN (\pp[24] [53] ), .A1 (n_0_39), .A2 (n_0_31));
NOR2_X1 i_0_292 (.ZN (\pp[24] [52] ), .A1 (n_0_39), .A2 (n_0_30));
NOR2_X1 i_0_291 (.ZN (\pp[24] [51] ), .A1 (n_0_39), .A2 (n_0_29));
NOR2_X1 i_0_290 (.ZN (\pp[24] [50] ), .A1 (n_0_39), .A2 (n_0_28));
NOR2_X1 i_0_289 (.ZN (\pp[24] [49] ), .A1 (n_0_39), .A2 (n_0_27));
NOR2_X1 i_0_288 (.ZN (\pp[24] [48] ), .A1 (n_0_39), .A2 (n_0_26));
NOR2_X1 i_0_287 (.ZN (\pp[24] [47] ), .A1 (n_0_39), .A2 (n_0_25));
NOR2_X1 i_0_286 (.ZN (\pp[24] [46] ), .A1 (n_0_39), .A2 (n_0_24));
NOR2_X1 i_0_285 (.ZN (\pp[24] [45] ), .A1 (n_0_39), .A2 (n_0_23));
NOR2_X1 i_0_284 (.ZN (\pp[24] [44] ), .A1 (n_0_39), .A2 (n_0_22));
NOR2_X1 i_0_283 (.ZN (\pp[24] [43] ), .A1 (n_0_39), .A2 (n_0_21));
NOR2_X1 i_0_282 (.ZN (\pp[24] [42] ), .A1 (n_0_39), .A2 (n_0_20));
NOR2_X1 i_0_281 (.ZN (\pp[24] [41] ), .A1 (n_0_39), .A2 (n_0_19));
NOR2_X1 i_0_280 (.ZN (\pp[24] [40] ), .A1 (n_0_39), .A2 (n_0_18));
NOR2_X1 i_0_279 (.ZN (\pp[24] [39] ), .A1 (n_0_39), .A2 (n_0_17));
NOR2_X1 i_0_278 (.ZN (\pp[24] [38] ), .A1 (n_0_39), .A2 (n_0_16));
NOR2_X1 i_0_277 (.ZN (\pp[24] [37] ), .A1 (n_0_39), .A2 (sgo__n50));
NOR2_X1 i_0_276 (.ZN (\pp[24] [36] ), .A1 (n_0_39), .A2 (sgo__n240));
NOR2_X1 i_0_275 (.ZN (\pp[24] [35] ), .A1 (n_0_39), .A2 (sgo__n106));
NOR2_X1 i_0_274 (.ZN (\pp[24] [34] ), .A1 (n_0_39), .A2 (sgo__n157));
NOR2_X1 i_0_273 (.ZN (\pp[24] [33] ), .A1 (n_0_39), .A2 (sgo__n133));
NOR2_X1 i_0_272 (.ZN (\pp[24] [32] ), .A1 (n_0_39), .A2 (sgo__n162));
NOR2_X1 i_0_271 (.ZN (\pp[24] [31] ), .A1 (n_0_39), .A2 (sgo__n74));
NOR2_X1 i_0_270 (.ZN (\pp[24] [30] ), .A1 (n_0_39), .A2 (sgo__n184));
NOR2_X1 i_0_269 (.ZN (\pp[24] [29] ), .A1 (n_0_39), .A2 (sgo__n172));
NOR2_X1 i_0_268 (.ZN (\pp[24] [28] ), .A1 (n_0_39), .A2 (sgo__n147));
NOR2_X1 i_0_267 (.ZN (\pp[24] [27] ), .A1 (n_0_39), .A2 (n_0_5));
NOR2_X1 i_0_266 (.ZN (\pp[24] [26] ), .A1 (n_0_39), .A2 (n_0_4));
NOR2_X1 i_0_265 (.ZN (\pp[24] [25] ), .A1 (n_0_39), .A2 (n_0_3));
NOR2_X1 i_0_264 (.ZN (\pp[24] [24] ), .A1 (n_0_39), .A2 (n_0_2));
INV_X4 i_0_263 (.ZN (n_0_39), .A (x[24]));
NOR2_X1 i_0_262 (.ZN (\pp[25] [63] ), .A1 (n_0_38), .A2 (n_0_33));
NOR2_X1 i_0_261 (.ZN (\pp[25] [55] ), .A1 (n_0_38), .A2 (n_0_32));
NOR2_X1 i_0_260 (.ZN (\pp[25] [54] ), .A1 (n_0_38), .A2 (n_0_31));
NOR2_X1 i_0_259 (.ZN (\pp[25] [53] ), .A1 (n_0_38), .A2 (n_0_30));
NOR2_X1 i_0_258 (.ZN (\pp[25] [52] ), .A1 (n_0_38), .A2 (n_0_29));
NOR2_X1 i_0_257 (.ZN (\pp[25] [51] ), .A1 (n_0_38), .A2 (n_0_28));
NOR2_X1 i_0_256 (.ZN (\pp[25] [50] ), .A1 (n_0_38), .A2 (n_0_27));
NOR2_X1 i_0_255 (.ZN (\pp[25] [49] ), .A1 (n_0_38), .A2 (n_0_26));
NOR2_X1 i_0_254 (.ZN (\pp[25] [48] ), .A1 (n_0_38), .A2 (n_0_25));
NOR2_X1 i_0_253 (.ZN (\pp[25] [47] ), .A1 (n_0_38), .A2 (n_0_24));
NOR2_X1 i_0_252 (.ZN (\pp[25] [46] ), .A1 (n_0_38), .A2 (n_0_23));
NOR2_X1 i_0_251 (.ZN (\pp[25] [45] ), .A1 (n_0_38), .A2 (n_0_22));
NOR2_X1 i_0_250 (.ZN (\pp[25] [44] ), .A1 (n_0_38), .A2 (n_0_21));
NOR2_X1 i_0_249 (.ZN (\pp[25] [43] ), .A1 (n_0_38), .A2 (n_0_20));
NOR2_X1 i_0_248 (.ZN (\pp[25] [42] ), .A1 (n_0_38), .A2 (n_0_19));
NOR2_X1 i_0_247 (.ZN (\pp[25] [41] ), .A1 (n_0_38), .A2 (n_0_18));
NOR2_X1 i_0_246 (.ZN (\pp[25] [40] ), .A1 (n_0_38), .A2 (n_0_17));
NOR2_X1 i_0_245 (.ZN (\pp[25] [39] ), .A1 (n_0_38), .A2 (n_0_16));
NOR2_X1 i_0_244 (.ZN (\pp[25] [38] ), .A1 (n_0_38), .A2 (sgo__n50));
NOR2_X1 i_0_243 (.ZN (\pp[25] [37] ), .A1 (n_0_38), .A2 (sgo__n240));
NOR2_X1 i_0_242 (.ZN (\pp[25] [36] ), .A1 (n_0_38), .A2 (sgo__n106));
NOR2_X1 i_0_241 (.ZN (\pp[25] [35] ), .A1 (n_0_38), .A2 (sgo__n157));
NOR2_X1 i_0_240 (.ZN (\pp[25] [34] ), .A1 (n_0_38), .A2 (sgo__n133));
NOR2_X1 i_0_239 (.ZN (\pp[25] [33] ), .A1 (n_0_38), .A2 (sgo__n162));
NOR2_X1 i_0_238 (.ZN (\pp[25] [32] ), .A1 (n_0_38), .A2 (sgo__n74));
NOR2_X1 i_0_237 (.ZN (\pp[25] [31] ), .A1 (n_0_38), .A2 (sgo__n184));
NOR2_X1 i_0_236 (.ZN (\pp[25] [30] ), .A1 (n_0_38), .A2 (sgo__n172));
NOR2_X1 i_0_235 (.ZN (\pp[25] [29] ), .A1 (n_0_38), .A2 (sgo__n147));
NOR2_X1 i_0_234 (.ZN (\pp[25] [28] ), .A1 (n_0_38), .A2 (n_0_5));
NOR2_X1 i_0_233 (.ZN (\pp[25] [27] ), .A1 (n_0_38), .A2 (slo___n701));
NOR2_X1 i_0_232 (.ZN (\pp[25] [26] ), .A1 (n_0_38), .A2 (n_0_3));
NOR2_X1 i_0_231 (.ZN (\pp[25] [25] ), .A1 (n_0_38), .A2 (n_0_2));
INV_X2 i_0_230 (.ZN (n_0_38), .A (x[25]));
NOR2_X1 i_0_229 (.ZN (\pp[26] [63] ), .A1 (n_0_37), .A2 (n_0_33));
NOR2_X1 i_0_228 (.ZN (\pp[26] [56] ), .A1 (n_0_37), .A2 (n_0_32));
NOR2_X1 i_0_227 (.ZN (\pp[26] [55] ), .A1 (n_0_37), .A2 (n_0_31));
NOR2_X1 i_0_226 (.ZN (\pp[26] [54] ), .A1 (n_0_37), .A2 (n_0_30));
NOR2_X1 i_0_225 (.ZN (\pp[26] [53] ), .A1 (n_0_37), .A2 (n_0_29));
NOR2_X1 i_0_224 (.ZN (\pp[26] [52] ), .A1 (n_0_37), .A2 (n_0_28));
NOR2_X1 i_0_223 (.ZN (\pp[26] [51] ), .A1 (n_0_37), .A2 (n_0_27));
NOR2_X1 i_0_222 (.ZN (\pp[26] [50] ), .A1 (n_0_37), .A2 (n_0_26));
NOR2_X1 i_0_221 (.ZN (\pp[26] [49] ), .A1 (n_0_37), .A2 (n_0_25));
NOR2_X1 i_0_220 (.ZN (\pp[26] [48] ), .A1 (n_0_37), .A2 (n_0_24));
NOR2_X1 i_0_219 (.ZN (\pp[26] [47] ), .A1 (n_0_37), .A2 (n_0_23));
NOR2_X1 i_0_218 (.ZN (\pp[26] [46] ), .A1 (n_0_37), .A2 (n_0_22));
NOR2_X1 i_0_217 (.ZN (\pp[26] [45] ), .A1 (n_0_37), .A2 (n_0_21));
NOR2_X1 i_0_216 (.ZN (\pp[26] [44] ), .A1 (n_0_37), .A2 (n_0_20));
NOR2_X1 i_0_215 (.ZN (\pp[26] [43] ), .A1 (n_0_37), .A2 (n_0_19));
NOR2_X1 i_0_214 (.ZN (\pp[26] [42] ), .A1 (n_0_37), .A2 (n_0_18));
NOR2_X1 i_0_213 (.ZN (\pp[26] [41] ), .A1 (n_0_37), .A2 (n_0_17));
NOR2_X1 i_0_212 (.ZN (\pp[26] [40] ), .A1 (n_0_37), .A2 (n_0_16));
NOR2_X1 i_0_211 (.ZN (\pp[26] [39] ), .A1 (n_0_37), .A2 (sgo__n50));
NOR2_X1 i_0_210 (.ZN (\pp[26] [38] ), .A1 (n_0_37), .A2 (sgo__n240));
NOR2_X1 i_0_209 (.ZN (\pp[26] [37] ), .A1 (n_0_37), .A2 (sgo__n106));
NOR2_X1 i_0_208 (.ZN (\pp[26] [36] ), .A1 (n_0_37), .A2 (sgo__n157));
NOR2_X1 i_0_207 (.ZN (\pp[26] [35] ), .A1 (n_0_37), .A2 (sgo__n133));
NOR2_X1 i_0_206 (.ZN (\pp[26] [34] ), .A1 (n_0_37), .A2 (sgo__n162));
NOR2_X1 i_0_205 (.ZN (\pp[26] [33] ), .A1 (n_0_37), .A2 (sgo__n74));
NOR2_X1 i_0_204 (.ZN (\pp[26] [32] ), .A1 (n_0_37), .A2 (sgo__n184));
NOR2_X1 i_0_203 (.ZN (\pp[26] [31] ), .A1 (n_0_37), .A2 (sgo__n172));
NOR2_X1 i_0_202 (.ZN (\pp[26] [30] ), .A1 (n_0_37), .A2 (sgo__n147));
NOR2_X1 i_0_201 (.ZN (\pp[26] [29] ), .A1 (n_0_37), .A2 (n_0_5));
NOR2_X1 i_0_200 (.ZN (\pp[26] [28] ), .A1 (n_0_37), .A2 (slo___n701));
NOR2_X1 i_0_199 (.ZN (\pp[26] [27] ), .A1 (n_0_37), .A2 (n_0_3));
NOR2_X1 i_0_198 (.ZN (\pp[26] [26] ), .A1 (n_0_37), .A2 (n_0_2));
INV_X2 i_0_197 (.ZN (n_0_37), .A (x[26]));
NOR2_X1 i_0_196 (.ZN (\pp[27] [63] ), .A1 (n_0_36), .A2 (n_0_33));
NOR2_X1 i_0_195 (.ZN (\pp[27] [57] ), .A1 (n_0_36), .A2 (n_0_32));
NOR2_X1 i_0_194 (.ZN (\pp[27] [56] ), .A1 (n_0_36), .A2 (n_0_31));
NOR2_X1 i_0_193 (.ZN (\pp[27] [55] ), .A1 (n_0_36), .A2 (n_0_30));
NOR2_X1 i_0_192 (.ZN (\pp[27] [54] ), .A1 (n_0_36), .A2 (n_0_29));
NOR2_X1 i_0_191 (.ZN (\pp[27] [53] ), .A1 (n_0_36), .A2 (n_0_28));
NOR2_X1 i_0_190 (.ZN (\pp[27] [52] ), .A1 (n_0_36), .A2 (n_0_27));
NOR2_X1 i_0_189 (.ZN (\pp[27] [51] ), .A1 (n_0_36), .A2 (n_0_26));
NOR2_X1 i_0_188 (.ZN (\pp[27] [50] ), .A1 (n_0_36), .A2 (n_0_25));
NOR2_X1 i_0_187 (.ZN (\pp[27] [49] ), .A1 (n_0_36), .A2 (n_0_24));
NOR2_X1 i_0_186 (.ZN (\pp[27] [48] ), .A1 (n_0_36), .A2 (n_0_23));
NOR2_X1 i_0_185 (.ZN (\pp[27] [47] ), .A1 (n_0_36), .A2 (n_0_22));
NOR2_X1 i_0_184 (.ZN (\pp[27] [46] ), .A1 (n_0_36), .A2 (n_0_21));
NOR2_X1 i_0_183 (.ZN (\pp[27] [45] ), .A1 (n_0_36), .A2 (n_0_20));
NOR2_X1 i_0_182 (.ZN (\pp[27] [44] ), .A1 (n_0_36), .A2 (n_0_19));
NOR2_X1 i_0_181 (.ZN (\pp[27] [43] ), .A1 (n_0_36), .A2 (n_0_18));
NOR2_X1 i_0_180 (.ZN (\pp[27] [42] ), .A1 (n_0_36), .A2 (n_0_17));
NOR2_X1 i_0_179 (.ZN (\pp[27] [41] ), .A1 (n_0_36), .A2 (n_0_16));
NOR2_X1 i_0_178 (.ZN (\pp[27] [40] ), .A1 (n_0_36), .A2 (sgo__n50));
NOR2_X1 i_0_177 (.ZN (\pp[27] [39] ), .A1 (n_0_36), .A2 (sgo__n240));
NOR2_X1 i_0_176 (.ZN (\pp[27] [38] ), .A1 (n_0_36), .A2 (sgo__n106));
NOR2_X1 i_0_175 (.ZN (\pp[27] [37] ), .A1 (n_0_36), .A2 (sgo__n157));
NOR2_X1 i_0_174 (.ZN (\pp[27] [36] ), .A1 (n_0_36), .A2 (sgo__n133));
NOR2_X1 i_0_173 (.ZN (\pp[27] [35] ), .A1 (n_0_36), .A2 (sgo__n162));
NOR2_X1 i_0_172 (.ZN (\pp[27] [34] ), .A1 (n_0_36), .A2 (sgo__n74));
NOR2_X1 i_0_171 (.ZN (\pp[27] [33] ), .A1 (n_0_36), .A2 (sgo__n184));
NOR2_X1 i_0_170 (.ZN (\pp[27] [32] ), .A1 (n_0_36), .A2 (sgo__n172));
NOR2_X1 i_0_169 (.ZN (\pp[27] [31] ), .A1 (n_0_36), .A2 (sgo__n147));
NOR2_X1 i_0_168 (.ZN (\pp[27] [30] ), .A1 (n_0_36), .A2 (n_0_5));
NOR2_X1 i_0_167 (.ZN (\pp[27] [29] ), .A1 (n_0_36), .A2 (slo___n701));
NOR2_X1 i_0_166 (.ZN (\pp[27] [28] ), .A1 (n_0_36), .A2 (n_0_3));
NOR2_X1 i_0_165 (.ZN (\pp[27] [27] ), .A1 (n_0_36), .A2 (n_0_2));
INV_X2 i_0_164 (.ZN (n_0_36), .A (x[27]));
NOR2_X1 i_0_163 (.ZN (\pp[28] [63] ), .A1 (n_0_35), .A2 (n_0_33));
NOR2_X1 i_0_162 (.ZN (\pp[28] [58] ), .A1 (n_0_35), .A2 (n_0_32));
NOR2_X1 i_0_161 (.ZN (\pp[28] [57] ), .A1 (n_0_35), .A2 (n_0_31));
NOR2_X1 i_0_160 (.ZN (\pp[28] [56] ), .A1 (n_0_35), .A2 (n_0_30));
NOR2_X1 i_0_159 (.ZN (\pp[28] [55] ), .A1 (n_0_35), .A2 (n_0_29));
NOR2_X1 i_0_158 (.ZN (\pp[28] [54] ), .A1 (n_0_35), .A2 (n_0_28));
NOR2_X1 i_0_157 (.ZN (\pp[28] [53] ), .A1 (n_0_35), .A2 (n_0_27));
NOR2_X1 i_0_156 (.ZN (\pp[28] [52] ), .A1 (n_0_35), .A2 (n_0_26));
NOR2_X1 i_0_155 (.ZN (\pp[28] [51] ), .A1 (n_0_35), .A2 (n_0_25));
NOR2_X1 i_0_154 (.ZN (\pp[28] [50] ), .A1 (n_0_35), .A2 (n_0_24));
NOR2_X1 i_0_153 (.ZN (\pp[28] [49] ), .A1 (n_0_35), .A2 (n_0_23));
NOR2_X1 i_0_152 (.ZN (\pp[28] [48] ), .A1 (n_0_35), .A2 (n_0_22));
NOR2_X1 i_0_151 (.ZN (\pp[28] [47] ), .A1 (n_0_35), .A2 (n_0_21));
NOR2_X1 i_0_150 (.ZN (\pp[28] [46] ), .A1 (n_0_35), .A2 (n_0_20));
NOR2_X1 i_0_149 (.ZN (\pp[28] [45] ), .A1 (n_0_35), .A2 (n_0_19));
NOR2_X1 i_0_148 (.ZN (\pp[28] [44] ), .A1 (n_0_35), .A2 (n_0_18));
NOR2_X1 i_0_147 (.ZN (\pp[28] [43] ), .A1 (n_0_35), .A2 (n_0_17));
NOR2_X1 i_0_146 (.ZN (\pp[28] [42] ), .A1 (n_0_35), .A2 (n_0_16));
NOR2_X1 i_0_145 (.ZN (\pp[28] [41] ), .A1 (n_0_35), .A2 (sgo__n50));
NOR2_X1 i_0_144 (.ZN (\pp[28] [40] ), .A1 (n_0_35), .A2 (sgo__n240));
NOR2_X1 i_0_143 (.ZN (\pp[28] [39] ), .A1 (n_0_35), .A2 (sgo__n106));
NOR2_X1 i_0_142 (.ZN (\pp[28] [38] ), .A1 (n_0_35), .A2 (sgo__n157));
NOR2_X1 i_0_141 (.ZN (\pp[28] [37] ), .A1 (n_0_35), .A2 (sgo__n133));
NOR2_X1 i_0_140 (.ZN (\pp[28] [36] ), .A1 (n_0_35), .A2 (sgo__n162));
NOR2_X1 i_0_139 (.ZN (\pp[28] [35] ), .A1 (n_0_35), .A2 (sgo__n74));
NOR2_X1 i_0_138 (.ZN (\pp[28] [34] ), .A1 (n_0_35), .A2 (sgo__n184));
NOR2_X1 i_0_137 (.ZN (\pp[28] [33] ), .A1 (n_0_35), .A2 (sgo__n172));
NOR2_X1 i_0_136 (.ZN (\pp[28] [32] ), .A1 (n_0_35), .A2 (sgo__n147));
NOR2_X1 i_0_135 (.ZN (\pp[28] [31] ), .A1 (n_0_35), .A2 (n_0_5));
NOR2_X1 i_0_134 (.ZN (\pp[28] [30] ), .A1 (n_0_35), .A2 (slo___n701));
NOR2_X1 i_0_133 (.ZN (\pp[28] [29] ), .A1 (n_0_35), .A2 (n_0_3));
NOR2_X1 i_0_132 (.ZN (\pp[28] [28] ), .A1 (n_0_35), .A2 (n_0_2));
INV_X2 i_0_131 (.ZN (n_0_35), .A (x[28]));
NOR2_X1 i_0_130 (.ZN (\pp[29] [63] ), .A1 (n_0_34), .A2 (n_0_33));
NOR2_X1 i_0_129 (.ZN (\pp[29] [59] ), .A1 (n_0_34), .A2 (n_0_32));
NOR2_X1 i_0_128 (.ZN (\pp[29] [58] ), .A1 (n_0_34), .A2 (n_0_31));
NOR2_X1 i_0_127 (.ZN (\pp[29] [57] ), .A1 (n_0_34), .A2 (n_0_30));
NOR2_X1 i_0_126 (.ZN (\pp[29] [56] ), .A1 (n_0_34), .A2 (n_0_29));
NOR2_X1 i_0_125 (.ZN (\pp[29] [55] ), .A1 (n_0_34), .A2 (n_0_28));
NOR2_X1 i_0_124 (.ZN (\pp[29] [54] ), .A1 (n_0_34), .A2 (n_0_27));
NOR2_X1 i_0_123 (.ZN (\pp[29] [53] ), .A1 (n_0_34), .A2 (n_0_26));
NOR2_X1 i_0_122 (.ZN (\pp[29] [52] ), .A1 (n_0_34), .A2 (n_0_25));
NOR2_X1 i_0_121 (.ZN (\pp[29] [51] ), .A1 (n_0_34), .A2 (n_0_24));
NOR2_X1 i_0_120 (.ZN (\pp[29] [50] ), .A1 (n_0_34), .A2 (n_0_23));
NOR2_X1 i_0_119 (.ZN (\pp[29] [49] ), .A1 (n_0_34), .A2 (n_0_22));
NOR2_X1 i_0_118 (.ZN (\pp[29] [48] ), .A1 (n_0_34), .A2 (n_0_21));
NOR2_X1 i_0_117 (.ZN (\pp[29] [47] ), .A1 (n_0_34), .A2 (n_0_20));
NOR2_X1 i_0_116 (.ZN (\pp[29] [46] ), .A1 (n_0_34), .A2 (n_0_19));
NOR2_X1 i_0_115 (.ZN (\pp[29] [45] ), .A1 (n_0_34), .A2 (n_0_18));
NOR2_X1 i_0_114 (.ZN (\pp[29] [44] ), .A1 (n_0_34), .A2 (n_0_17));
NOR2_X1 i_0_113 (.ZN (\pp[29] [43] ), .A1 (n_0_34), .A2 (n_0_16));
NOR2_X1 i_0_112 (.ZN (\pp[29] [42] ), .A1 (n_0_34), .A2 (sgo__n50));
NOR2_X1 i_0_111 (.ZN (\pp[29] [41] ), .A1 (n_0_34), .A2 (sgo__n240));
NOR2_X1 i_0_110 (.ZN (\pp[29] [40] ), .A1 (n_0_34), .A2 (sgo__n106));
NOR2_X1 i_0_109 (.ZN (\pp[29] [39] ), .A1 (n_0_34), .A2 (sgo__n157));
NOR2_X1 i_0_108 (.ZN (\pp[29] [38] ), .A1 (n_0_34), .A2 (sgo__n133));
NOR2_X1 i_0_107 (.ZN (\pp[29] [37] ), .A1 (n_0_34), .A2 (sgo__n162));
NOR2_X1 i_0_106 (.ZN (\pp[29] [36] ), .A1 (n_0_34), .A2 (sgo__n74));
NOR2_X1 i_0_105 (.ZN (\pp[29] [35] ), .A1 (n_0_34), .A2 (sgo__n184));
NOR2_X1 i_0_104 (.ZN (\pp[29] [34] ), .A1 (n_0_34), .A2 (sgo__n172));
NOR2_X1 i_0_103 (.ZN (\pp[29] [33] ), .A1 (n_0_34), .A2 (sgo__n147));
NOR2_X1 i_0_102 (.ZN (\pp[29] [32] ), .A1 (n_0_34), .A2 (n_0_5));
NOR2_X1 i_0_101 (.ZN (\pp[29] [31] ), .A1 (n_0_34), .A2 (slo___n701));
NOR2_X1 i_0_100 (.ZN (\pp[29] [30] ), .A1 (n_0_34), .A2 (n_0_3));
NOR2_X1 i_0_99 (.ZN (\pp[29] [29] ), .A1 (n_0_34), .A2 (n_0_2));
INV_X2 i_0_98 (.ZN (n_0_34), .A (x[29]));
NOR2_X1 i_0_97 (.ZN (\pp[30] [63] ), .A1 (n_0_1), .A2 (n_0_33));
INV_X2 i_0_96 (.ZN (n_0_33), .A (y[31]));
NOR2_X1 i_0_95 (.ZN (\pp[30] [60] ), .A1 (n_0_1), .A2 (n_0_32));
INV_X2 i_0_94 (.ZN (n_0_32), .A (y[30]));
NOR2_X1 i_0_93 (.ZN (\pp[30] [59] ), .A1 (n_0_1), .A2 (n_0_31));
INV_X2 i_0_92 (.ZN (n_0_31), .A (y[29]));
NOR2_X1 i_0_91 (.ZN (\pp[30] [58] ), .A1 (n_0_1), .A2 (n_0_30));
INV_X2 i_0_90 (.ZN (n_0_30), .A (y[28]));
NOR2_X1 i_0_89 (.ZN (\pp[30] [57] ), .A1 (n_0_1), .A2 (n_0_29));
INV_X2 i_0_88 (.ZN (n_0_29), .A (y[27]));
NOR2_X1 i_0_87 (.ZN (\pp[30] [56] ), .A1 (n_0_1), .A2 (n_0_28));
INV_X2 i_0_86 (.ZN (n_0_28), .A (y[26]));
NOR2_X1 i_0_85 (.ZN (\pp[30] [55] ), .A1 (n_0_1), .A2 (n_0_27));
INV_X2 i_0_84 (.ZN (n_0_27), .A (y[25]));
NOR2_X1 i_0_83 (.ZN (\pp[30] [54] ), .A1 (n_0_1), .A2 (n_0_26));
INV_X2 i_0_82 (.ZN (n_0_26), .A (y[24]));
NOR2_X1 i_0_81 (.ZN (\pp[30] [53] ), .A1 (n_0_1), .A2 (n_0_25));
INV_X2 i_0_80 (.ZN (n_0_25), .A (y[23]));
NOR2_X1 i_0_79 (.ZN (\pp[30] [52] ), .A1 (n_0_1), .A2 (n_0_24));
INV_X2 i_0_78 (.ZN (n_0_24), .A (y[22]));
NOR2_X1 i_0_77 (.ZN (\pp[30] [51] ), .A1 (n_0_1), .A2 (n_0_23));
INV_X2 i_0_76 (.ZN (n_0_23), .A (y[21]));
NOR2_X1 i_0_75 (.ZN (\pp[30] [50] ), .A1 (n_0_1), .A2 (n_0_22));
INV_X2 i_0_74 (.ZN (n_0_22), .A (y[20]));
NOR2_X1 i_0_73 (.ZN (\pp[30] [49] ), .A1 (n_0_1), .A2 (n_0_21));
INV_X4 i_0_72 (.ZN (n_0_21), .A (y[19]));
NOR2_X1 i_0_71 (.ZN (\pp[30] [48] ), .A1 (n_0_1), .A2 (n_0_20));
INV_X4 i_0_70 (.ZN (n_0_20), .A (y[18]));
NOR2_X1 i_0_69 (.ZN (\pp[30] [47] ), .A1 (n_0_1), .A2 (n_0_19));
INV_X8 i_0_68 (.ZN (n_0_19), .A (y[17]));
NOR2_X1 i_0_67 (.ZN (\pp[30] [46] ), .A1 (n_0_1), .A2 (n_0_18));
INV_X8 i_0_66 (.ZN (n_0_18), .A (y[16]));
NOR2_X1 i_0_65 (.ZN (\pp[30] [45] ), .A1 (n_0_1), .A2 (n_0_17));
INV_X8 i_0_64 (.ZN (n_0_17), .A (y[15]));
NOR2_X1 i_0_63 (.ZN (\pp[30] [44] ), .A1 (n_0_1), .A2 (n_0_16));
INV_X8 i_0_62 (.ZN (n_0_16), .A (y[14]));
NOR2_X1 i_0_61 (.ZN (\pp[30] [43] ), .A1 (n_0_1), .A2 (sgo__n50));
INV_X8 i_0_60 (.ZN (n_0_15), .A (y[13]));
NOR2_X1 i_0_59 (.ZN (\pp[30] [42] ), .A1 (n_0_1), .A2 (sgo__n240));
INV_X16 i_0_58 (.ZN (n_0_14), .A (y[12]));
NOR2_X1 i_0_57 (.ZN (\pp[30] [41] ), .A1 (n_0_1), .A2 (sgo__n106));
NOR2_X1 i_0_55 (.ZN (\pp[30] [40] ), .A1 (n_0_1), .A2 (sgo__n157));
NOR2_X1 i_0_53 (.ZN (\pp[30] [39] ), .A1 (n_0_1), .A2 (sgo__n133));
NOR2_X1 i_0_51 (.ZN (\pp[30] [38] ), .A1 (n_0_1), .A2 (sgo__n162));
NOR2_X1 i_0_49 (.ZN (\pp[30] [37] ), .A1 (n_0_1), .A2 (sgo__n74));
NOR2_X1 i_0_47 (.ZN (\pp[30] [36] ), .A1 (n_0_1), .A2 (sgo__n184));
NOR2_X1 i_0_45 (.ZN (\pp[30] [35] ), .A1 (n_0_1), .A2 (sgo__n172));
NOR2_X1 i_0_43 (.ZN (\pp[30] [34] ), .A1 (n_0_1), .A2 (sgo__n147));
NOR2_X1 i_0_41 (.ZN (\pp[30] [33] ), .A1 (n_0_1), .A2 (n_0_5));
NOR2_X1 i_0_39 (.ZN (\pp[30] [32] ), .A1 (n_0_1), .A2 (slo___n701));
NOR2_X1 i_0_37 (.ZN (\pp[30] [31] ), .A1 (n_0_1), .A2 (n_0_3));
INV_X8 i_0_36 (.ZN (n_0_3), .A (y[1]));
NOR2_X1 i_0_35 (.ZN (\pp[30] [30] ), .A1 (n_0_1), .A2 (n_0_2));
INV_X8 i_0_34 (.ZN (n_0_2), .A (y[0]));
INV_X2 i_0_33 (.ZN (n_0_1), .A (x[30]));
NOR2_X1 i_0_32 (.ZN (\pp[31] [63] ), .A1 (n_0_0), .A2 (y[31]));
NOR2_X1 i_0_31 (.ZN (\pp[31] [61] ), .A1 (n_0_0), .A2 (y[30]));
NOR2_X1 i_0_30 (.ZN (\pp[31] [60] ), .A1 (n_0_0), .A2 (y[29]));
NOR2_X1 i_0_29 (.ZN (\pp[31] [59] ), .A1 (n_0_0), .A2 (y[28]));
NOR2_X1 i_0_28 (.ZN (\pp[31] [58] ), .A1 (n_0_0), .A2 (y[27]));
NOR2_X1 i_0_27 (.ZN (\pp[31] [57] ), .A1 (n_0_0), .A2 (y[26]));
NOR2_X1 i_0_26 (.ZN (\pp[31] [56] ), .A1 (n_0_0), .A2 (y[25]));
NOR2_X1 i_0_25 (.ZN (\pp[31] [55] ), .A1 (n_0_0), .A2 (y[24]));
NOR2_X1 i_0_24 (.ZN (\pp[31] [54] ), .A1 (n_0_0), .A2 (y[23]));
NOR2_X1 i_0_23 (.ZN (\pp[31] [53] ), .A1 (n_0_0), .A2 (y[22]));
NOR2_X1 i_0_22 (.ZN (\pp[31] [52] ), .A1 (n_0_0), .A2 (y[21]));
NOR2_X1 i_0_21 (.ZN (\pp[31] [51] ), .A1 (n_0_0), .A2 (y[20]));
NOR2_X1 i_0_20 (.ZN (\pp[31] [50] ), .A1 (n_0_0), .A2 (y[19]));
NOR2_X1 i_0_19 (.ZN (\pp[31] [49] ), .A1 (n_0_0), .A2 (y[18]));
NOR2_X1 i_0_18 (.ZN (\pp[31] [48] ), .A1 (n_0_0), .A2 (y[17]));
NOR2_X1 i_0_17 (.ZN (\pp[31] [47] ), .A1 (n_0_0), .A2 (y[16]));
NOR2_X1 i_0_16 (.ZN (\pp[31] [46] ), .A1 (n_0_0), .A2 (y[15]));
NOR2_X1 i_0_15 (.ZN (\pp[31] [45] ), .A1 (n_0_0), .A2 (y[14]));
NOR2_X1 i_0_14 (.ZN (\pp[31] [44] ), .A1 (n_0_0), .A2 (y[13]));
NOR2_X2 i_0_13 (.ZN (\pp[31] [43] ), .A1 (n_0_0), .A2 (y[12]));
NOR2_X2 i_0_12 (.ZN (\pp[31] [42] ), .A1 (n_0_0), .A2 (y[11]));
NOR2_X1 i_0_11 (.ZN (\pp[31] [41] ), .A1 (n_0_0), .A2 (y[10]));
NOR2_X1 i_0_10 (.ZN (\pp[31] [40] ), .A1 (n_0_0), .A2 (y[9]));
NOR2_X1 i_0_9 (.ZN (\pp[31] [39] ), .A1 (n_0_0), .A2 (y[8]));
NOR2_X1 i_0_8 (.ZN (\pp[31] [38] ), .A1 (n_0_0), .A2 (y[7]));
NOR2_X2 i_0_7 (.ZN (\pp[31] [37] ), .A1 (n_0_0), .A2 (y[6]));
NOR2_X1 i_0_6 (.ZN (\pp[31] [36] ), .A1 (n_0_0), .A2 (y[5]));
NOR2_X1 i_0_5 (.ZN (\pp[31] [35] ), .A1 (n_0_0), .A2 (y[4]));
NOR2_X1 i_0_4 (.ZN (\pp[31] [34] ), .A1 (n_0_0), .A2 (y[3]));
NOR2_X1 i_0_3 (.ZN (\pp[31] [33] ), .A1 (n_0_0), .A2 (y[2]));
NOR2_X1 i_0_2 (.ZN (\pp[31] [32] ), .A1 (n_0_0), .A2 (y[1]));
NOR2_X1 i_0_1 (.ZN (\pp[31] [31] ), .A1 (n_0_0), .A2 (y[0]));
INV_X4 i_0_0 (.ZN (n_0_0), .A (x[31]));
BUF_X16 sgo__c150 (.Z (sgo__n150), .A (n_0_60));
BUF_X2 sgo__c160 (.Z (sgo__n157), .A (n_0_12));
BUF_X8 sgo__c168 (.Z (sgo__n162), .A (n_0_10));
BUF_X8 sgo__c176 (.Z (sgo__n167), .A (n_0_61));
BUF_X16 sgo__c184 (.Z (sgo__n172), .A (n_0_7));
BUF_X4 sgo__c192 (.Z (sgo__n177), .A (n_0_11));
BUF_X8 sgo__c202 (.Z (sgo__n184), .A (n_0_8));
BUF_X8 sgo__c225 (.Z (sgo__n205), .A (sgo__n149));
CLKBUF_X3 sgo__c265 (.Z (sgo__n240), .A (n_0_14));
BUF_X8 sgo__c302 (.Z (sgo__n272), .A (n_0_55));
BUF_X16 sgo__c334 (.Z (sgo__n301), .A (n_0_63));
NOR2_X2 slo__sro_c534 (.ZN (\pp[9] [11] ), .A1 (n_0_4), .A2 (n_0_54));
BUF_X8 slo__c459 (.Z (slo__n415), .A (n_0_61));
BUF_X8 sgo__c354 (.Z (sgo__n315), .A (n_0_59));
BUF_X4 sgo__L1_c31 (.Z (sgo__n31), .A (n_0_3));
BUF_X1 sgo__L1_c34 (.Z (sgo__n34), .A (n_0_3));
BUF_X8 sgo__L1_c39 (.Z (sgo__n39), .A (n_0_2));
CLKBUF_X2 slo___L1_c591 (.Z (slo___n553), .A (n_0_58));
INV_X4 slo__c618 (.ZN (slo__n580), .A (y[4]));
NAND2_X4 slo__sro_c638 (.ZN (slo__sro_n602), .A1 (x[2]), .A2 (y[8]));
BUF_X2 sgo__L1_c46 (.Z (sgo__n46), .A (n_0_15));
BUF_X1 sgo__L1_c48 (.Z (sgo__n48), .A (n_0_15));
BUF_X1 sgo__L1_c50 (.Z (sgo__n50), .A (n_0_15));
INV_X4 slo__sro_c639 (.ZN (\pp[2] [10] ), .A (slo__sro_n602));
BUF_X4 drc_ipo_c947 (.Z (drc_ipo_n910), .A (n_0_43));
BUF_X2 sgo__L1_c66 (.Z (sgo__n66), .A (n_0_4));
BUF_X1 sgo__L4_c69 (.Z (sgo__n69), .A (sgo__n66));
BUF_X1 sgo__L4_c74 (.Z (sgo__n74), .A (n_0_9));
BUF_X2 sgo__L1_c106 (.Z (sgo__n106), .A (n_0_13));
BUF_X4 drc_ipo_c948 (.Z (drc_ipo_n911), .A (n_0_42));
NOR2_X4 slo__sro_c1055 (.ZN (\pp[11] [12] ), .A1 (sgo__n31), .A2 (n_0_52));
BUF_X1 sgo__L1_c133 (.Z (sgo__n133), .A (sgo__n177));
BUF_X1 sgo__L1_c140 (.Z (sgo__n140), .A (sgo__n240));
BUF_X1 sgo__L1_c147 (.Z (sgo__n147), .A (n_0_6));
BUF_X8 sgo__L1_c149 (.Z (sgo__n149), .A (slo__n580));

endmodule //products

module mulTree (x, y, out);

output [63:0] out;
input [31:0] x;
input [31:0] y;
wire \pp[0][63] ;
wire \pp[0][30] ;
wire \pp[0][29] ;
wire \pp[0][28] ;
wire \pp[0][27] ;
wire \pp[0][26] ;
wire \pp[0][25] ;
wire \pp[0][24] ;
wire \pp[0][23] ;
wire \pp[0][22] ;
wire \pp[0][21] ;
wire \pp[0][20] ;
wire \pp[0][19] ;
wire \pp[0][18] ;
wire \pp[0][17] ;
wire \pp[0][16] ;
wire \pp[0][15] ;
wire \pp[0][14] ;
wire \pp[0][13] ;
wire \pp[0][12] ;
wire \pp[0][11] ;
wire \pp[0][10] ;
wire \pp[0][9] ;
wire \pp[0][8] ;
wire \pp[0][7] ;
wire \pp[0][6] ;
wire \pp[0][5] ;
wire \pp[0][4] ;
wire \pp[0][3] ;
wire \pp[0][2] ;
wire \pp[0][1] ;
wire \pp[1][63] ;
wire \pp[1][31] ;
wire \pp[1][30] ;
wire \pp[1][29] ;
wire \pp[1][28] ;
wire \pp[1][27] ;
wire \pp[1][26] ;
wire \pp[1][25] ;
wire \pp[1][24] ;
wire \pp[1][23] ;
wire \pp[1][22] ;
wire \pp[1][21] ;
wire \pp[1][20] ;
wire \pp[1][19] ;
wire \pp[1][18] ;
wire \pp[1][17] ;
wire \pp[1][16] ;
wire \pp[1][15] ;
wire \pp[1][14] ;
wire \pp[1][13] ;
wire \pp[1][12] ;
wire \pp[1][11] ;
wire \pp[1][10] ;
wire \pp[1][9] ;
wire \pp[1][8] ;
wire \pp[1][7] ;
wire \pp[1][6] ;
wire \pp[1][5] ;
wire \pp[1][4] ;
wire \pp[1][3] ;
wire \pp[1][2] ;
wire \pp[1][1] ;
wire \pp[2][63] ;
wire \pp[2][32] ;
wire \pp[2][31] ;
wire \pp[2][30] ;
wire \pp[2][29] ;
wire \pp[2][28] ;
wire \pp[2][27] ;
wire \pp[2][26] ;
wire \pp[2][25] ;
wire \pp[2][24] ;
wire \pp[2][23] ;
wire \pp[2][22] ;
wire \pp[2][21] ;
wire \pp[2][20] ;
wire \pp[2][19] ;
wire \pp[2][18] ;
wire \pp[2][17] ;
wire \pp[2][16] ;
wire \pp[2][15] ;
wire \pp[2][14] ;
wire \pp[2][13] ;
wire \pp[2][12] ;
wire \pp[2][11] ;
wire \pp[2][10] ;
wire \pp[2][9] ;
wire \pp[2][8] ;
wire \pp[2][7] ;
wire \pp[2][6] ;
wire \pp[2][5] ;
wire \pp[2][4] ;
wire \pp[2][3] ;
wire \pp[2][2] ;
wire \pp[3][63] ;
wire \pp[3][33] ;
wire \pp[3][32] ;
wire \pp[3][31] ;
wire \pp[3][30] ;
wire \pp[3][29] ;
wire \pp[3][28] ;
wire \pp[3][27] ;
wire \pp[3][26] ;
wire \pp[3][25] ;
wire \pp[3][24] ;
wire \pp[3][23] ;
wire \pp[3][22] ;
wire \pp[3][21] ;
wire \pp[3][20] ;
wire \pp[3][19] ;
wire \pp[3][18] ;
wire \pp[3][17] ;
wire \pp[3][16] ;
wire \pp[3][15] ;
wire \pp[3][14] ;
wire \pp[3][13] ;
wire \pp[3][12] ;
wire \pp[3][11] ;
wire \pp[3][10] ;
wire \pp[3][9] ;
wire \pp[3][8] ;
wire \pp[3][7] ;
wire \pp[3][6] ;
wire \pp[3][5] ;
wire \pp[3][4] ;
wire \pp[3][3] ;
wire \pp[4][63] ;
wire \pp[4][34] ;
wire \pp[4][33] ;
wire \pp[4][32] ;
wire \pp[4][31] ;
wire \pp[4][30] ;
wire \pp[4][29] ;
wire \pp[4][28] ;
wire \pp[4][27] ;
wire \pp[4][26] ;
wire \pp[4][25] ;
wire \pp[4][24] ;
wire \pp[4][23] ;
wire \pp[4][22] ;
wire \pp[4][21] ;
wire \pp[4][20] ;
wire \pp[4][19] ;
wire \pp[4][18] ;
wire \pp[4][17] ;
wire \pp[4][16] ;
wire \pp[4][15] ;
wire \pp[4][14] ;
wire \pp[4][13] ;
wire \pp[4][12] ;
wire \pp[4][11] ;
wire \pp[4][10] ;
wire \pp[4][9] ;
wire \pp[4][8] ;
wire \pp[4][7] ;
wire \pp[4][6] ;
wire \pp[4][5] ;
wire \pp[4][4] ;
wire \pp[5][63] ;
wire \pp[5][35] ;
wire \pp[5][34] ;
wire \pp[5][33] ;
wire \pp[5][32] ;
wire \pp[5][31] ;
wire \pp[5][30] ;
wire \pp[5][29] ;
wire \pp[5][28] ;
wire \pp[5][27] ;
wire \pp[5][26] ;
wire \pp[5][25] ;
wire \pp[5][24] ;
wire \pp[5][23] ;
wire \pp[5][22] ;
wire \pp[5][21] ;
wire \pp[5][20] ;
wire \pp[5][19] ;
wire \pp[5][18] ;
wire \pp[5][17] ;
wire \pp[5][16] ;
wire \pp[5][15] ;
wire \pp[5][14] ;
wire \pp[5][13] ;
wire \pp[5][12] ;
wire \pp[5][11] ;
wire \pp[5][10] ;
wire \pp[5][9] ;
wire \pp[5][8] ;
wire \pp[5][7] ;
wire \pp[5][6] ;
wire \pp[5][5] ;
wire \pp[6][63] ;
wire \pp[6][36] ;
wire \pp[6][35] ;
wire \pp[6][34] ;
wire \pp[6][33] ;
wire \pp[6][32] ;
wire \pp[6][31] ;
wire \pp[6][30] ;
wire \pp[6][29] ;
wire \pp[6][28] ;
wire \pp[6][27] ;
wire \pp[6][26] ;
wire \pp[6][25] ;
wire \pp[6][24] ;
wire \pp[6][23] ;
wire \pp[6][22] ;
wire \pp[6][21] ;
wire \pp[6][20] ;
wire \pp[6][19] ;
wire \pp[6][18] ;
wire \pp[6][17] ;
wire \pp[6][16] ;
wire \pp[6][15] ;
wire \pp[6][14] ;
wire \pp[6][13] ;
wire \pp[6][12] ;
wire \pp[6][11] ;
wire \pp[6][10] ;
wire \pp[6][9] ;
wire \pp[6][8] ;
wire \pp[6][7] ;
wire \pp[6][6] ;
wire \pp[7][63] ;
wire \pp[7][37] ;
wire \pp[7][36] ;
wire \pp[7][35] ;
wire \pp[7][34] ;
wire \pp[7][33] ;
wire \pp[7][32] ;
wire \pp[7][31] ;
wire \pp[7][30] ;
wire \pp[7][29] ;
wire \pp[7][28] ;
wire \pp[7][27] ;
wire \pp[7][26] ;
wire \pp[7][25] ;
wire \pp[7][24] ;
wire \pp[7][23] ;
wire \pp[7][22] ;
wire \pp[7][21] ;
wire \pp[7][20] ;
wire \pp[7][19] ;
wire \pp[7][18] ;
wire \pp[7][17] ;
wire \pp[7][16] ;
wire \pp[7][15] ;
wire \pp[7][14] ;
wire \pp[7][13] ;
wire \pp[7][12] ;
wire \pp[7][11] ;
wire \pp[7][10] ;
wire \pp[7][9] ;
wire \pp[7][8] ;
wire \pp[7][7] ;
wire \pp[8][63] ;
wire \pp[8][38] ;
wire \pp[8][37] ;
wire \pp[8][36] ;
wire \pp[8][35] ;
wire \pp[8][34] ;
wire \pp[8][33] ;
wire \pp[8][32] ;
wire \pp[8][31] ;
wire \pp[8][30] ;
wire \pp[8][29] ;
wire \pp[8][28] ;
wire \pp[8][27] ;
wire \pp[8][26] ;
wire \pp[8][25] ;
wire \pp[8][24] ;
wire \pp[8][23] ;
wire \pp[8][22] ;
wire \pp[8][21] ;
wire \pp[8][20] ;
wire \pp[8][19] ;
wire \pp[8][18] ;
wire \pp[8][17] ;
wire \pp[8][16] ;
wire \pp[8][15] ;
wire \pp[8][14] ;
wire \pp[8][13] ;
wire \pp[8][12] ;
wire \pp[8][11] ;
wire \pp[8][10] ;
wire \pp[8][9] ;
wire \pp[8][8] ;
wire \pp[9][63] ;
wire \pp[9][39] ;
wire \pp[9][38] ;
wire \pp[9][37] ;
wire \pp[9][36] ;
wire \pp[9][35] ;
wire \pp[9][34] ;
wire \pp[9][33] ;
wire \pp[9][32] ;
wire \pp[9][31] ;
wire \pp[9][30] ;
wire \pp[9][29] ;
wire \pp[9][28] ;
wire \pp[9][27] ;
wire \pp[9][26] ;
wire \pp[9][25] ;
wire \pp[9][24] ;
wire \pp[9][23] ;
wire \pp[9][22] ;
wire \pp[9][21] ;
wire \pp[9][20] ;
wire \pp[9][19] ;
wire \pp[9][18] ;
wire \pp[9][17] ;
wire \pp[9][16] ;
wire \pp[9][15] ;
wire \pp[9][14] ;
wire \pp[9][13] ;
wire \pp[9][12] ;
wire \pp[9][11] ;
wire \pp[9][10] ;
wire \pp[9][9] ;
wire \pp[10][63] ;
wire \pp[10][40] ;
wire \pp[10][39] ;
wire \pp[10][38] ;
wire \pp[10][37] ;
wire \pp[10][36] ;
wire \pp[10][35] ;
wire \pp[10][34] ;
wire \pp[10][33] ;
wire \pp[10][32] ;
wire \pp[10][31] ;
wire \pp[10][30] ;
wire \pp[10][29] ;
wire \pp[10][28] ;
wire \pp[10][27] ;
wire \pp[10][26] ;
wire \pp[10][25] ;
wire \pp[10][24] ;
wire \pp[10][23] ;
wire \pp[10][22] ;
wire \pp[10][21] ;
wire \pp[10][20] ;
wire \pp[10][19] ;
wire \pp[10][18] ;
wire \pp[10][17] ;
wire \pp[10][16] ;
wire \pp[10][15] ;
wire \pp[10][14] ;
wire \pp[10][13] ;
wire \pp[10][12] ;
wire \pp[10][11] ;
wire \pp[10][10] ;
wire \pp[11][63] ;
wire \pp[11][41] ;
wire \pp[11][40] ;
wire \pp[11][39] ;
wire \pp[11][38] ;
wire \pp[11][37] ;
wire \pp[11][36] ;
wire \pp[11][35] ;
wire \pp[11][34] ;
wire \pp[11][33] ;
wire \pp[11][32] ;
wire \pp[11][31] ;
wire \pp[11][30] ;
wire \pp[11][29] ;
wire \pp[11][28] ;
wire \pp[11][27] ;
wire \pp[11][26] ;
wire \pp[11][25] ;
wire \pp[11][24] ;
wire \pp[11][23] ;
wire \pp[11][22] ;
wire \pp[11][21] ;
wire \pp[11][20] ;
wire \pp[11][19] ;
wire \pp[11][18] ;
wire \pp[11][17] ;
wire \pp[11][16] ;
wire \pp[11][15] ;
wire \pp[11][14] ;
wire \pp[11][13] ;
wire \pp[11][12] ;
wire \pp[11][11] ;
wire \sums[4][63] ;
wire \sums[4][44] ;
wire \sums[4][43] ;
wire \sums[4][42] ;
wire \sums[4][41] ;
wire \sums[4][40] ;
wire \sums[4][39] ;
wire \sums[4][38] ;
wire \sums[4][37] ;
wire \sums[4][36] ;
wire \sums[4][35] ;
wire \sums[4][34] ;
wire \sums[4][33] ;
wire \sums[4][32] ;
wire \sums[4][31] ;
wire \sums[4][30] ;
wire \sums[4][29] ;
wire \sums[4][28] ;
wire \sums[4][27] ;
wire \sums[4][26] ;
wire \sums[4][25] ;
wire \sums[4][24] ;
wire \sums[4][23] ;
wire \sums[4][22] ;
wire \sums[4][21] ;
wire \sums[4][20] ;
wire \sums[4][19] ;
wire \sums[4][18] ;
wire \sums[4][17] ;
wire \sums[4][16] ;
wire \sums[4][15] ;
wire \sums[4][14] ;
wire \sums[4][13] ;
wire \sums[4][12] ;
wire \pp[12][62] ;
wire \pp[12][42] ;
wire \pp[12][41] ;
wire \pp[12][40] ;
wire \pp[12][39] ;
wire \pp[12][38] ;
wire \pp[12][37] ;
wire \pp[12][36] ;
wire \pp[12][35] ;
wire \pp[12][34] ;
wire \pp[12][33] ;
wire \pp[12][32] ;
wire \pp[12][31] ;
wire \pp[12][30] ;
wire \pp[12][29] ;
wire \pp[12][28] ;
wire \pp[12][27] ;
wire \pp[12][26] ;
wire \pp[12][25] ;
wire \pp[12][24] ;
wire \pp[12][23] ;
wire \pp[12][22] ;
wire \pp[12][21] ;
wire \pp[12][20] ;
wire \pp[12][19] ;
wire \pp[12][18] ;
wire \pp[12][17] ;
wire \pp[12][16] ;
wire \pp[12][15] ;
wire \pp[12][14] ;
wire \pp[12][13] ;
wire \pp[13][62] ;
wire \pp[13][43] ;
wire \pp[13][42] ;
wire \pp[13][41] ;
wire \pp[13][40] ;
wire \pp[13][39] ;
wire \pp[13][38] ;
wire \pp[13][37] ;
wire \pp[13][36] ;
wire \pp[13][35] ;
wire \pp[13][34] ;
wire \pp[13][33] ;
wire \pp[13][32] ;
wire \pp[13][31] ;
wire \pp[13][30] ;
wire \pp[13][29] ;
wire \pp[13][28] ;
wire \pp[13][27] ;
wire \pp[13][26] ;
wire \pp[13][25] ;
wire \pp[13][24] ;
wire \pp[13][23] ;
wire \pp[13][22] ;
wire \pp[13][21] ;
wire \pp[13][20] ;
wire \pp[13][19] ;
wire \pp[13][18] ;
wire \pp[13][17] ;
wire \pp[13][16] ;
wire \pp[13][15] ;
wire \pp[13][14] ;
wire \pp[13][13] ;
wire \pp[14][62] ;
wire \pp[14][44] ;
wire \pp[14][43] ;
wire \pp[14][42] ;
wire \pp[14][41] ;
wire \pp[14][40] ;
wire \pp[14][39] ;
wire \pp[14][38] ;
wire \pp[14][37] ;
wire \pp[14][36] ;
wire \pp[14][35] ;
wire \pp[14][34] ;
wire \pp[14][33] ;
wire \pp[14][32] ;
wire \pp[14][31] ;
wire \pp[14][30] ;
wire \pp[14][29] ;
wire \pp[14][28] ;
wire \pp[14][27] ;
wire \pp[14][26] ;
wire \pp[14][25] ;
wire \pp[14][24] ;
wire \pp[14][23] ;
wire \pp[14][22] ;
wire \pp[14][21] ;
wire \pp[14][20] ;
wire \pp[14][19] ;
wire \pp[14][18] ;
wire \pp[14][17] ;
wire \pp[14][16] ;
wire \pp[14][15] ;
wire \pp[14][14] ;
wire \pp[15][62] ;
wire \pp[15][45] ;
wire \pp[15][44] ;
wire \pp[15][43] ;
wire \pp[15][42] ;
wire \pp[15][41] ;
wire \pp[15][40] ;
wire \pp[15][39] ;
wire \pp[15][38] ;
wire \pp[15][37] ;
wire \pp[15][36] ;
wire \pp[15][35] ;
wire \pp[15][34] ;
wire \pp[15][33] ;
wire \pp[15][32] ;
wire \pp[15][31] ;
wire \pp[15][30] ;
wire \pp[15][29] ;
wire \pp[15][28] ;
wire \pp[15][27] ;
wire \pp[15][26] ;
wire \pp[15][25] ;
wire \pp[15][24] ;
wire \pp[15][23] ;
wire \pp[15][22] ;
wire \pp[15][21] ;
wire \pp[15][20] ;
wire \pp[15][19] ;
wire \pp[15][18] ;
wire \pp[15][17] ;
wire \pp[15][16] ;
wire \pp[15][15] ;
wire \pp[16][62] ;
wire \pp[16][46] ;
wire \pp[16][45] ;
wire \pp[16][44] ;
wire \pp[16][43] ;
wire \pp[16][42] ;
wire \pp[16][41] ;
wire \pp[16][40] ;
wire \pp[16][39] ;
wire \pp[16][38] ;
wire \pp[16][37] ;
wire \pp[16][36] ;
wire \pp[16][35] ;
wire \pp[16][34] ;
wire \pp[16][33] ;
wire \pp[16][32] ;
wire \pp[16][31] ;
wire \pp[16][30] ;
wire \pp[16][29] ;
wire \pp[16][28] ;
wire \pp[16][27] ;
wire \pp[16][26] ;
wire \pp[16][25] ;
wire \pp[16][24] ;
wire \pp[16][23] ;
wire \pp[16][22] ;
wire \pp[16][21] ;
wire \pp[16][20] ;
wire \pp[16][19] ;
wire \pp[16][18] ;
wire \pp[16][17] ;
wire \pp[16][16] ;
wire \pp[17][62] ;
wire \pp[17][47] ;
wire \pp[17][46] ;
wire \pp[17][45] ;
wire \pp[17][44] ;
wire \pp[17][43] ;
wire \pp[17][42] ;
wire \pp[17][41] ;
wire \pp[17][40] ;
wire \pp[17][39] ;
wire \pp[17][38] ;
wire \pp[17][37] ;
wire \pp[17][36] ;
wire \pp[17][35] ;
wire \pp[17][34] ;
wire \pp[17][33] ;
wire \pp[17][32] ;
wire \pp[17][31] ;
wire \pp[17][30] ;
wire \pp[17][29] ;
wire \pp[17][28] ;
wire \pp[17][27] ;
wire \pp[17][26] ;
wire \pp[17][25] ;
wire \pp[17][24] ;
wire \pp[17][23] ;
wire \pp[17][22] ;
wire \pp[17][21] ;
wire \pp[17][20] ;
wire \pp[17][19] ;
wire \pp[17][18] ;
wire \pp[17][17] ;
wire \pp[18][63] ;
wire \pp[18][48] ;
wire \pp[18][47] ;
wire \pp[18][46] ;
wire \pp[18][45] ;
wire \pp[18][44] ;
wire \pp[18][43] ;
wire \pp[18][42] ;
wire \pp[18][41] ;
wire \pp[18][40] ;
wire \pp[18][39] ;
wire \pp[18][38] ;
wire \pp[18][37] ;
wire \pp[18][36] ;
wire \pp[18][35] ;
wire \pp[18][34] ;
wire \pp[18][33] ;
wire \pp[18][32] ;
wire \pp[18][31] ;
wire \pp[18][30] ;
wire \pp[18][29] ;
wire \pp[18][28] ;
wire \pp[18][27] ;
wire \pp[18][26] ;
wire \pp[18][25] ;
wire \pp[18][24] ;
wire \pp[18][23] ;
wire \pp[18][22] ;
wire \pp[18][21] ;
wire \pp[18][20] ;
wire \pp[18][19] ;
wire \pp[18][18] ;
wire \pp[19][63] ;
wire \pp[19][49] ;
wire \pp[19][48] ;
wire \pp[19][47] ;
wire \pp[19][46] ;
wire \pp[19][45] ;
wire \pp[19][44] ;
wire \pp[19][43] ;
wire \pp[19][42] ;
wire \pp[19][41] ;
wire \pp[19][40] ;
wire \pp[19][39] ;
wire \pp[19][38] ;
wire \pp[19][37] ;
wire \pp[19][36] ;
wire \pp[19][35] ;
wire \pp[19][34] ;
wire \pp[19][33] ;
wire \pp[19][32] ;
wire \pp[19][31] ;
wire \pp[19][30] ;
wire \pp[19][29] ;
wire \pp[19][28] ;
wire \pp[19][27] ;
wire \pp[19][26] ;
wire \pp[19][25] ;
wire \pp[19][24] ;
wire \pp[19][23] ;
wire \pp[19][22] ;
wire \pp[19][21] ;
wire \pp[19][20] ;
wire \pp[19][19] ;
wire \pp[20][63] ;
wire \pp[20][50] ;
wire \pp[20][49] ;
wire \pp[20][48] ;
wire \pp[20][47] ;
wire \pp[20][46] ;
wire \pp[20][45] ;
wire \pp[20][44] ;
wire \pp[20][43] ;
wire \pp[20][42] ;
wire \pp[20][41] ;
wire \pp[20][40] ;
wire \pp[20][39] ;
wire \pp[20][38] ;
wire \pp[20][37] ;
wire \pp[20][36] ;
wire \pp[20][35] ;
wire \pp[20][34] ;
wire \pp[20][33] ;
wire \pp[20][32] ;
wire \pp[20][31] ;
wire \pp[20][30] ;
wire \pp[20][29] ;
wire \pp[20][28] ;
wire \pp[20][27] ;
wire \pp[20][26] ;
wire \pp[20][25] ;
wire \pp[20][24] ;
wire \pp[20][23] ;
wire \pp[20][22] ;
wire \pp[20][21] ;
wire \pp[20][20] ;
wire \pp[21][63] ;
wire \pp[21][51] ;
wire \pp[21][50] ;
wire \pp[21][49] ;
wire \pp[21][48] ;
wire \pp[21][47] ;
wire \pp[21][46] ;
wire \pp[21][45] ;
wire \pp[21][44] ;
wire \pp[21][43] ;
wire \pp[21][42] ;
wire \pp[21][41] ;
wire \pp[21][40] ;
wire \pp[21][39] ;
wire \pp[21][38] ;
wire \pp[21][37] ;
wire \pp[21][36] ;
wire \pp[21][35] ;
wire \pp[21][34] ;
wire \pp[21][33] ;
wire \pp[21][32] ;
wire \pp[21][31] ;
wire \pp[21][30] ;
wire \pp[21][29] ;
wire \pp[21][28] ;
wire \pp[21][27] ;
wire \pp[21][26] ;
wire \pp[21][25] ;
wire \pp[21][24] ;
wire \pp[21][23] ;
wire \pp[21][22] ;
wire \pp[21][21] ;
wire \pp[22][63] ;
wire \pp[22][52] ;
wire \pp[22][51] ;
wire \pp[22][50] ;
wire \pp[22][49] ;
wire \pp[22][48] ;
wire \pp[22][47] ;
wire \pp[22][46] ;
wire \pp[22][45] ;
wire \pp[22][44] ;
wire \pp[22][43] ;
wire \pp[22][42] ;
wire \pp[22][41] ;
wire \pp[22][40] ;
wire \pp[22][39] ;
wire \pp[22][38] ;
wire \pp[22][37] ;
wire \pp[22][36] ;
wire \pp[22][35] ;
wire \pp[22][34] ;
wire \pp[22][33] ;
wire \pp[22][32] ;
wire \pp[22][31] ;
wire \pp[22][30] ;
wire \pp[22][29] ;
wire \pp[22][28] ;
wire \pp[22][27] ;
wire \pp[22][26] ;
wire \pp[22][25] ;
wire \pp[22][24] ;
wire \pp[22][23] ;
wire \pp[22][22] ;
wire \pp[23][63] ;
wire \pp[23][53] ;
wire \pp[23][52] ;
wire \pp[23][51] ;
wire \pp[23][50] ;
wire \pp[23][49] ;
wire \pp[23][48] ;
wire \pp[23][47] ;
wire \pp[23][46] ;
wire \pp[23][45] ;
wire \pp[23][44] ;
wire \pp[23][43] ;
wire \pp[23][42] ;
wire \pp[23][41] ;
wire \pp[23][40] ;
wire \pp[23][39] ;
wire \pp[23][38] ;
wire \pp[23][37] ;
wire \pp[23][36] ;
wire \pp[23][35] ;
wire \pp[23][34] ;
wire \pp[23][33] ;
wire \pp[23][32] ;
wire \pp[23][31] ;
wire \pp[23][30] ;
wire \pp[23][29] ;
wire \pp[23][28] ;
wire \pp[23][27] ;
wire \pp[23][26] ;
wire \pp[23][25] ;
wire \pp[23][24] ;
wire \pp[23][23] ;
wire \pp[24][63] ;
wire \pp[24][54] ;
wire \pp[24][53] ;
wire \pp[24][52] ;
wire \pp[24][51] ;
wire \pp[24][50] ;
wire \pp[24][49] ;
wire \pp[24][48] ;
wire \pp[24][47] ;
wire \pp[24][46] ;
wire \pp[24][45] ;
wire \pp[24][44] ;
wire \pp[24][43] ;
wire \pp[24][42] ;
wire \pp[24][41] ;
wire \pp[24][40] ;
wire \pp[24][39] ;
wire \pp[24][38] ;
wire \pp[24][37] ;
wire \pp[24][36] ;
wire \pp[24][35] ;
wire \pp[24][34] ;
wire \pp[24][33] ;
wire \pp[24][32] ;
wire \pp[24][31] ;
wire \pp[24][30] ;
wire \pp[24][29] ;
wire \pp[24][28] ;
wire \pp[24][27] ;
wire \pp[24][26] ;
wire \pp[24][25] ;
wire \pp[24][24] ;
wire \pp[25][63] ;
wire \pp[25][55] ;
wire \pp[25][54] ;
wire \pp[25][53] ;
wire \pp[25][52] ;
wire \pp[25][51] ;
wire \pp[25][50] ;
wire \pp[25][49] ;
wire \pp[25][48] ;
wire \pp[25][47] ;
wire \pp[25][46] ;
wire \pp[25][45] ;
wire \pp[25][44] ;
wire \pp[25][43] ;
wire \pp[25][42] ;
wire \pp[25][41] ;
wire \pp[25][40] ;
wire \pp[25][39] ;
wire \pp[25][38] ;
wire \pp[25][37] ;
wire \pp[25][36] ;
wire \pp[25][35] ;
wire \pp[25][34] ;
wire \pp[25][33] ;
wire \pp[25][32] ;
wire \pp[25][31] ;
wire \pp[25][30] ;
wire \pp[25][29] ;
wire \pp[25][28] ;
wire \pp[25][27] ;
wire \pp[25][26] ;
wire \pp[25][25] ;
wire \pp[26][63] ;
wire \pp[26][56] ;
wire \pp[26][55] ;
wire \pp[26][54] ;
wire \pp[26][53] ;
wire \pp[26][52] ;
wire \pp[26][51] ;
wire \pp[26][50] ;
wire \pp[26][49] ;
wire \pp[26][48] ;
wire \pp[26][47] ;
wire \pp[26][46] ;
wire \pp[26][45] ;
wire \pp[26][44] ;
wire \pp[26][43] ;
wire \pp[26][42] ;
wire \pp[26][41] ;
wire \pp[26][40] ;
wire \pp[26][39] ;
wire \pp[26][38] ;
wire \pp[26][37] ;
wire \pp[26][36] ;
wire \pp[26][35] ;
wire \pp[26][34] ;
wire \pp[26][33] ;
wire \pp[26][32] ;
wire \pp[26][31] ;
wire \pp[26][30] ;
wire \pp[26][29] ;
wire \pp[26][28] ;
wire \pp[26][27] ;
wire \pp[26][26] ;
wire \pp[27][58] ;
wire \pp[27][57] ;
wire \pp[27][56] ;
wire \pp[27][55] ;
wire \pp[27][54] ;
wire \pp[27][53] ;
wire \pp[27][52] ;
wire \pp[27][51] ;
wire \pp[27][50] ;
wire \pp[27][49] ;
wire \pp[27][48] ;
wire \pp[27][47] ;
wire \pp[27][46] ;
wire \pp[27][45] ;
wire \pp[27][44] ;
wire \pp[27][43] ;
wire \pp[27][42] ;
wire \pp[27][41] ;
wire \pp[27][40] ;
wire \pp[27][39] ;
wire \pp[27][38] ;
wire \pp[27][37] ;
wire \pp[27][36] ;
wire \pp[27][35] ;
wire \pp[27][34] ;
wire \pp[27][33] ;
wire \pp[27][32] ;
wire \pp[27][31] ;
wire \pp[27][30] ;
wire \pp[27][29] ;
wire \pp[27][28] ;
wire \pp[27][27] ;
wire \pp[28][63] ;
wire \pp[28][58] ;
wire \pp[28][57] ;
wire \pp[28][56] ;
wire \pp[28][55] ;
wire \pp[28][54] ;
wire \pp[28][53] ;
wire \pp[28][52] ;
wire \pp[28][51] ;
wire \pp[28][50] ;
wire \pp[28][49] ;
wire \pp[28][48] ;
wire \pp[28][47] ;
wire \pp[28][46] ;
wire \pp[28][45] ;
wire \pp[28][44] ;
wire \pp[28][43] ;
wire \pp[28][42] ;
wire \pp[28][41] ;
wire \pp[28][40] ;
wire \pp[28][39] ;
wire \pp[28][38] ;
wire \pp[28][37] ;
wire \pp[28][36] ;
wire \pp[28][35] ;
wire \pp[28][34] ;
wire \pp[28][33] ;
wire \pp[28][32] ;
wire \pp[28][31] ;
wire \pp[28][30] ;
wire \pp[28][29] ;
wire \pp[28][28] ;
wire \pp[29][63] ;
wire \pp[29][59] ;
wire \pp[29][58] ;
wire \pp[29][57] ;
wire \pp[29][56] ;
wire \pp[29][55] ;
wire \pp[29][54] ;
wire \pp[29][53] ;
wire \pp[29][52] ;
wire \pp[29][51] ;
wire \pp[29][50] ;
wire \pp[29][49] ;
wire \pp[29][48] ;
wire \pp[29][47] ;
wire \pp[29][46] ;
wire \pp[29][45] ;
wire \pp[29][44] ;
wire \pp[29][43] ;
wire \pp[29][42] ;
wire \pp[29][41] ;
wire \pp[29][40] ;
wire \pp[29][39] ;
wire \pp[29][38] ;
wire \pp[29][37] ;
wire \pp[29][36] ;
wire \pp[29][35] ;
wire \pp[29][34] ;
wire \pp[29][33] ;
wire \pp[29][32] ;
wire \pp[29][31] ;
wire \pp[29][30] ;
wire \pp[29][29] ;
wire \pp[30][63] ;
wire \pp[30][60] ;
wire \pp[30][59] ;
wire \pp[30][58] ;
wire \pp[30][57] ;
wire \pp[30][56] ;
wire \pp[30][55] ;
wire \pp[30][54] ;
wire \pp[30][53] ;
wire \pp[30][52] ;
wire \pp[30][51] ;
wire \pp[30][50] ;
wire \pp[30][49] ;
wire \pp[30][48] ;
wire \pp[30][47] ;
wire \pp[30][46] ;
wire \pp[30][45] ;
wire \pp[30][44] ;
wire \pp[30][43] ;
wire \pp[30][42] ;
wire \pp[30][41] ;
wire \pp[30][40] ;
wire \pp[30][39] ;
wire \pp[30][38] ;
wire \pp[30][37] ;
wire \pp[30][36] ;
wire \pp[30][35] ;
wire \pp[30][34] ;
wire \pp[30][33] ;
wire \pp[30][32] ;
wire \pp[30][31] ;
wire \pp[30][30] ;
wire \pp[31][63] ;
wire \pp[31][61] ;
wire \pp[31][60] ;
wire \pp[31][59] ;
wire \pp[31][58] ;
wire \pp[31][57] ;
wire \pp[31][56] ;
wire \pp[31][55] ;
wire \pp[31][54] ;
wire \pp[31][53] ;
wire \pp[31][52] ;
wire \pp[31][51] ;
wire \pp[31][50] ;
wire \pp[31][49] ;
wire \pp[31][48] ;
wire \pp[31][47] ;
wire \pp[31][46] ;
wire \pp[31][45] ;
wire \pp[31][44] ;
wire \pp[31][43] ;
wire \pp[31][42] ;
wire \pp[31][41] ;
wire \pp[31][40] ;
wire \pp[31][39] ;
wire \pp[31][38] ;
wire \pp[31][37] ;
wire \pp[31][36] ;
wire \pp[31][35] ;
wire \pp[31][34] ;
wire \pp[31][33] ;
wire \pp[31][32] ;
wire \pp[31][31] ;
wire \couts[13][63] ;
wire \couts[13][49] ;
wire \couts[13][48] ;
wire \couts[13][47] ;
wire \couts[13][46] ;
wire \couts[13][45] ;
wire \couts[13][44] ;
wire \couts[13][43] ;
wire \couts[13][42] ;
wire \couts[13][41] ;
wire \couts[13][40] ;
wire \couts[13][39] ;
wire \couts[13][38] ;
wire \couts[13][37] ;
wire \couts[13][36] ;
wire \couts[13][35] ;
wire \couts[13][34] ;
wire \couts[13][33] ;
wire \couts[13][32] ;
wire \couts[13][31] ;
wire \couts[13][30] ;
wire \couts[13][29] ;
wire \couts[13][28] ;
wire \couts[13][27] ;
wire \couts[13][26] ;
wire \couts[13][25] ;
wire \couts[13][24] ;
wire \couts[13][23] ;
wire \couts[13][22] ;
wire \couts[13][21] ;
wire \couts[13][20] ;
wire \couts[13][19] ;
wire \couts[13][18] ;
wire \couts[13][17] ;
wire \couts[13][16] ;
wire \sums[13][63] ;
wire \sums[13][48] ;
wire \sums[13][47] ;
wire \sums[13][46] ;
wire \sums[13][45] ;
wire \sums[13][44] ;
wire \sums[13][43] ;
wire \sums[13][42] ;
wire \sums[13][41] ;
wire \sums[13][40] ;
wire \sums[13][39] ;
wire \sums[13][38] ;
wire \sums[13][37] ;
wire \sums[13][36] ;
wire \sums[13][35] ;
wire \sums[13][34] ;
wire \sums[13][33] ;
wire \sums[13][32] ;
wire \sums[13][31] ;
wire \sums[13][30] ;
wire \sums[13][29] ;
wire \sums[13][28] ;
wire \sums[13][27] ;
wire \sums[13][26] ;
wire \sums[13][25] ;
wire \sums[13][24] ;
wire \sums[13][23] ;
wire \sums[13][22] ;
wire \sums[13][21] ;
wire \sums[13][20] ;
wire \sums[13][19] ;
wire \sums[13][18] ;
wire \sums[13][17] ;
wire \sums[13][16] ;
wire \sums[13][15] ;
wire \sums[13][14] ;
wire \couts[5][63] ;
wire \couts[5][48] ;
wire \couts[5][47] ;
wire \couts[5][46] ;
wire \couts[5][45] ;
wire \couts[5][44] ;
wire \couts[5][43] ;
wire \couts[5][42] ;
wire \couts[5][41] ;
wire \couts[5][40] ;
wire \couts[5][39] ;
wire \couts[5][38] ;
wire \couts[5][37] ;
wire \couts[5][36] ;
wire \couts[5][35] ;
wire \couts[5][34] ;
wire \couts[5][33] ;
wire \couts[5][32] ;
wire \couts[5][31] ;
wire \couts[5][30] ;
wire \couts[5][29] ;
wire \couts[5][28] ;
wire \couts[5][27] ;
wire \couts[5][26] ;
wire \couts[5][25] ;
wire \couts[5][24] ;
wire \couts[5][23] ;
wire \couts[5][22] ;
wire \couts[5][21] ;
wire \couts[5][20] ;
wire \couts[5][19] ;
wire \couts[5][18] ;
wire \couts[5][17] ;
wire \sums[5][63] ;
wire \sums[5][47] ;
wire \sums[5][46] ;
wire \sums[5][45] ;
wire \sums[5][44] ;
wire \sums[5][43] ;
wire \sums[5][42] ;
wire \sums[5][41] ;
wire \sums[5][40] ;
wire \sums[5][39] ;
wire \sums[5][38] ;
wire \sums[5][37] ;
wire \sums[5][36] ;
wire \sums[5][35] ;
wire \sums[5][34] ;
wire \sums[5][33] ;
wire \sums[5][32] ;
wire \sums[5][31] ;
wire \sums[5][30] ;
wire \sums[5][29] ;
wire \sums[5][28] ;
wire \sums[5][27] ;
wire \sums[5][26] ;
wire \sums[5][25] ;
wire \sums[5][24] ;
wire \sums[5][23] ;
wire \sums[5][22] ;
wire \sums[5][21] ;
wire \sums[5][20] ;
wire \sums[5][19] ;
wire \sums[5][18] ;
wire \sums[5][17] ;
wire \sums[5][16] ;
wire \couts[4][63] ;
wire \couts[4][45] ;
wire \couts[4][44] ;
wire \couts[4][43] ;
wire \couts[4][42] ;
wire \couts[4][41] ;
wire \couts[4][40] ;
wire \couts[4][39] ;
wire \couts[4][38] ;
wire \couts[4][37] ;
wire \couts[4][36] ;
wire \couts[4][35] ;
wire \couts[4][34] ;
wire \couts[4][33] ;
wire \couts[4][32] ;
wire \couts[4][31] ;
wire \couts[4][30] ;
wire \couts[4][29] ;
wire \couts[4][28] ;
wire \couts[4][27] ;
wire \couts[4][26] ;
wire \couts[4][25] ;
wire \couts[4][24] ;
wire \couts[4][23] ;
wire \couts[4][22] ;
wire \couts[4][21] ;
wire \couts[4][20] ;
wire \couts[4][19] ;
wire \couts[4][18] ;
wire \couts[4][17] ;
wire \couts[4][16] ;
wire \couts[4][15] ;
wire \couts[2][63] ;
wire \couts[2][39] ;
wire \couts[2][38] ;
wire \couts[2][37] ;
wire \couts[2][36] ;
wire \couts[2][35] ;
wire \couts[2][34] ;
wire \couts[2][33] ;
wire \couts[2][32] ;
wire \couts[2][31] ;
wire \couts[2][30] ;
wire \couts[2][29] ;
wire \couts[2][28] ;
wire \couts[2][27] ;
wire \couts[2][26] ;
wire \couts[2][25] ;
wire \couts[2][24] ;
wire \couts[2][23] ;
wire \couts[2][22] ;
wire \couts[2][21] ;
wire \couts[2][20] ;
wire \couts[2][19] ;
wire \couts[2][18] ;
wire \couts[2][17] ;
wire \couts[2][16] ;
wire \couts[2][15] ;
wire \couts[2][14] ;
wire \couts[2][13] ;
wire \couts[2][12] ;
wire \couts[2][11] ;
wire \couts[2][10] ;
wire \couts[2][9] ;
wire \couts[2][8] ;
wire \sums[2][63] ;
wire \sums[2][38] ;
wire \sums[2][37] ;
wire \sums[2][36] ;
wire \sums[2][35] ;
wire \sums[2][34] ;
wire \sums[2][33] ;
wire \sums[2][32] ;
wire \sums[2][31] ;
wire \sums[2][30] ;
wire \sums[2][29] ;
wire \sums[2][28] ;
wire \sums[2][27] ;
wire \sums[2][26] ;
wire \sums[2][25] ;
wire \sums[2][24] ;
wire \sums[2][23] ;
wire \sums[2][22] ;
wire \sums[2][21] ;
wire \sums[2][20] ;
wire \sums[2][19] ;
wire \sums[2][18] ;
wire \sums[2][17] ;
wire \sums[2][16] ;
wire \sums[2][15] ;
wire \sums[2][14] ;
wire \sums[2][13] ;
wire \sums[2][12] ;
wire \sums[2][11] ;
wire \sums[2][10] ;
wire \sums[2][9] ;
wire \sums[2][8] ;
wire \sums[2][7] ;
wire \sums[18][63] ;
wire \sums[18][62] ;
wire \sums[18][61] ;
wire \sums[18][60] ;
wire \sums[18][59] ;
wire \sums[18][58] ;
wire \sums[18][57] ;
wire \sums[18][56] ;
wire \sums[18][55] ;
wire \sums[18][54] ;
wire \sums[18][53] ;
wire \sums[18][52] ;
wire \sums[18][51] ;
wire \sums[18][50] ;
wire \sums[18][49] ;
wire \sums[18][48] ;
wire \sums[18][47] ;
wire \sums[18][46] ;
wire \sums[18][45] ;
wire \sums[18][44] ;
wire \sums[18][43] ;
wire \sums[18][42] ;
wire \sums[18][41] ;
wire \sums[18][40] ;
wire \sums[18][39] ;
wire \sums[18][38] ;
wire \sums[18][37] ;
wire \sums[18][36] ;
wire \sums[18][35] ;
wire \sums[18][34] ;
wire \sums[18][33] ;
wire \sums[18][32] ;
wire \sums[18][31] ;
wire \sums[18][30] ;
wire \sums[18][29] ;
wire \sums[18][28] ;
wire \sums[18][27] ;
wire \sums[18][26] ;
wire \sums[18][25] ;
wire \sums[18][24] ;
wire \sums[18][23] ;
wire \sums[18][22] ;
wire \sums[18][21] ;
wire \sums[18][20] ;
wire \sums[18][19] ;
wire \sums[18][18] ;
wire \sums[18][17] ;
wire \sums[18][16] ;
wire \sums[18][15] ;
wire \sums[18][14] ;
wire \sums[18][13] ;
wire \sums[18][12] ;
wire \sums[18][11] ;
wire \sums[18][10] ;
wire \sums[18][9] ;
wire \sums[18][8] ;
wire \sums[18][7] ;
wire \couts[11][63] ;
wire \couts[11][62] ;
wire \couts[11][61] ;
wire \couts[11][60] ;
wire \couts[11][59] ;
wire \couts[11][58] ;
wire \couts[11][57] ;
wire \couts[11][56] ;
wire \couts[11][55] ;
wire \couts[11][54] ;
wire \couts[11][53] ;
wire \couts[11][52] ;
wire \couts[11][51] ;
wire \couts[11][50] ;
wire \couts[11][49] ;
wire \couts[11][48] ;
wire \couts[11][47] ;
wire \couts[11][46] ;
wire \couts[11][45] ;
wire \couts[11][44] ;
wire \couts[11][43] ;
wire \couts[11][42] ;
wire \couts[11][41] ;
wire \couts[11][40] ;
wire \couts[11][39] ;
wire \couts[11][38] ;
wire \couts[11][37] ;
wire \couts[11][36] ;
wire \couts[11][35] ;
wire \couts[11][34] ;
wire \couts[11][33] ;
wire \couts[11][32] ;
wire \couts[11][31] ;
wire \couts[11][30] ;
wire \couts[11][29] ;
wire \couts[11][28] ;
wire \couts[11][27] ;
wire \couts[11][26] ;
wire \couts[11][25] ;
wire \couts[11][24] ;
wire \couts[11][23] ;
wire \couts[11][22] ;
wire \couts[11][21] ;
wire \couts[11][20] ;
wire \couts[11][19] ;
wire \couts[11][18] ;
wire \couts[11][17] ;
wire \couts[11][16] ;
wire \couts[11][15] ;
wire \couts[11][14] ;
wire \couts[11][13] ;
wire \couts[11][12] ;
wire \couts[11][11] ;
wire \couts[11][10] ;
wire \couts[11][9] ;
wire \sums[11][63] ;
wire \sums[11][62] ;
wire \sums[11][61] ;
wire \sums[11][60] ;
wire \sums[11][59] ;
wire \sums[11][58] ;
wire \sums[11][57] ;
wire \sums[11][56] ;
wire \sums[11][55] ;
wire \sums[11][54] ;
wire \sums[11][53] ;
wire \sums[11][52] ;
wire \sums[11][51] ;
wire \sums[11][50] ;
wire \sums[11][49] ;
wire \sums[11][48] ;
wire \sums[11][47] ;
wire \sums[11][46] ;
wire \sums[11][45] ;
wire \sums[11][44] ;
wire \sums[11][43] ;
wire \sums[11][42] ;
wire \sums[11][41] ;
wire \sums[11][40] ;
wire \sums[11][39] ;
wire \sums[11][38] ;
wire \sums[11][37] ;
wire \sums[11][36] ;
wire \sums[11][35] ;
wire \sums[11][34] ;
wire \sums[11][33] ;
wire \sums[11][32] ;
wire \sums[11][31] ;
wire \sums[11][30] ;
wire \sums[11][29] ;
wire \sums[11][28] ;
wire \sums[11][27] ;
wire \sums[11][26] ;
wire \sums[11][25] ;
wire \sums[11][24] ;
wire \sums[11][23] ;
wire \sums[11][22] ;
wire \sums[11][21] ;
wire \sums[11][20] ;
wire \sums[11][19] ;
wire \sums[11][18] ;
wire \sums[11][17] ;
wire \sums[11][16] ;
wire \sums[11][15] ;
wire \sums[11][14] ;
wire \sums[11][13] ;
wire \sums[11][12] ;
wire \sums[11][11] ;
wire \sums[11][10] ;
wire \sums[11][9] ;
wire \sums[11][8] ;
wire \sums[11][7] ;
wire \sums[11][6] ;
wire \couts[12][63] ;
wire \couts[12][45] ;
wire \couts[12][44] ;
wire \couts[12][43] ;
wire \couts[12][42] ;
wire \couts[12][41] ;
wire \couts[12][40] ;
wire \couts[12][39] ;
wire \couts[12][38] ;
wire \couts[12][37] ;
wire \couts[12][36] ;
wire \couts[12][35] ;
wire \couts[12][34] ;
wire \couts[12][33] ;
wire \couts[12][32] ;
wire \couts[12][31] ;
wire \couts[12][30] ;
wire \couts[12][29] ;
wire \couts[12][28] ;
wire \couts[12][27] ;
wire \couts[12][26] ;
wire \couts[12][25] ;
wire \couts[12][24] ;
wire \couts[12][23] ;
wire \couts[12][22] ;
wire \couts[12][21] ;
wire \couts[12][20] ;
wire \couts[12][19] ;
wire \couts[12][18] ;
wire \couts[12][17] ;
wire \couts[12][16] ;
wire \couts[12][15] ;
wire \couts[12][14] ;
wire \couts[12][13] ;
wire \couts[12][12] ;
wire \sums[12][63] ;
wire \sums[12][44] ;
wire \sums[12][43] ;
wire \sums[12][42] ;
wire \sums[12][41] ;
wire \sums[12][40] ;
wire \sums[12][39] ;
wire \sums[12][38] ;
wire \sums[12][37] ;
wire \sums[12][36] ;
wire \sums[12][35] ;
wire \sums[12][34] ;
wire \sums[12][33] ;
wire \sums[12][32] ;
wire \sums[12][31] ;
wire \sums[12][30] ;
wire \sums[12][29] ;
wire \sums[12][28] ;
wire \sums[12][27] ;
wire \sums[12][26] ;
wire \sums[12][25] ;
wire \sums[12][24] ;
wire \sums[12][23] ;
wire \sums[12][22] ;
wire \sums[12][21] ;
wire \sums[12][20] ;
wire \sums[12][19] ;
wire \sums[12][18] ;
wire \sums[12][17] ;
wire \sums[12][16] ;
wire \sums[12][15] ;
wire \sums[12][14] ;
wire \sums[12][13] ;
wire \sums[12][12] ;
wire \sums[12][11] ;
wire \couts[3][63] ;
wire \couts[3][42] ;
wire \couts[3][41] ;
wire \couts[3][40] ;
wire \couts[3][39] ;
wire \couts[3][38] ;
wire \couts[3][37] ;
wire \couts[3][36] ;
wire \couts[3][35] ;
wire \couts[3][34] ;
wire \couts[3][33] ;
wire \couts[3][32] ;
wire \couts[3][31] ;
wire \couts[3][30] ;
wire \couts[3][29] ;
wire \couts[3][28] ;
wire \couts[3][27] ;
wire \couts[3][26] ;
wire \couts[3][25] ;
wire \couts[3][24] ;
wire \couts[3][23] ;
wire \couts[3][22] ;
wire \couts[3][21] ;
wire \couts[3][20] ;
wire \couts[3][19] ;
wire \couts[3][18] ;
wire \couts[3][17] ;
wire \couts[3][16] ;
wire \couts[3][15] ;
wire \couts[3][14] ;
wire \couts[3][13] ;
wire \couts[3][12] ;
wire \couts[3][11] ;
wire \sums[3][63] ;
wire \sums[3][41] ;
wire \sums[3][40] ;
wire \sums[3][39] ;
wire \sums[3][38] ;
wire \sums[3][37] ;
wire \sums[3][36] ;
wire \sums[3][35] ;
wire \sums[3][34] ;
wire \sums[3][33] ;
wire \sums[3][32] ;
wire \sums[3][31] ;
wire \sums[3][30] ;
wire \sums[3][29] ;
wire \sums[3][28] ;
wire \sums[3][27] ;
wire \sums[3][26] ;
wire \sums[3][25] ;
wire \sums[3][24] ;
wire \sums[3][23] ;
wire \sums[3][22] ;
wire \sums[3][21] ;
wire \sums[3][20] ;
wire \sums[3][19] ;
wire \sums[3][18] ;
wire \sums[3][17] ;
wire \sums[3][16] ;
wire \sums[3][15] ;
wire \sums[3][14] ;
wire \sums[3][13] ;
wire \sums[3][12] ;
wire \sums[3][11] ;
wire \sums[3][10] ;
wire \couts[18][63] ;
wire \couts[18][62] ;
wire \couts[18][61] ;
wire \couts[18][60] ;
wire \couts[18][59] ;
wire \couts[18][58] ;
wire \couts[18][57] ;
wire \couts[18][56] ;
wire \couts[18][55] ;
wire \couts[18][54] ;
wire \couts[18][53] ;
wire \couts[18][52] ;
wire \couts[18][51] ;
wire \couts[18][50] ;
wire \couts[18][49] ;
wire \couts[18][48] ;
wire \couts[18][47] ;
wire \couts[18][46] ;
wire \couts[18][45] ;
wire \couts[18][44] ;
wire \couts[18][43] ;
wire \couts[18][42] ;
wire \couts[18][41] ;
wire \couts[18][40] ;
wire \couts[18][39] ;
wire \couts[18][38] ;
wire \couts[18][37] ;
wire \couts[18][36] ;
wire \couts[18][35] ;
wire \couts[18][34] ;
wire \couts[18][33] ;
wire \couts[18][32] ;
wire \couts[18][31] ;
wire \couts[18][30] ;
wire \couts[18][29] ;
wire \couts[18][28] ;
wire \couts[18][27] ;
wire \couts[18][26] ;
wire \couts[18][25] ;
wire \couts[18][24] ;
wire \couts[18][23] ;
wire \couts[18][22] ;
wire \couts[18][21] ;
wire \couts[18][20] ;
wire \couts[18][19] ;
wire \couts[18][18] ;
wire \couts[18][17] ;
wire \couts[18][16] ;
wire \couts[18][15] ;
wire \couts[18][14] ;
wire \couts[18][13] ;
wire \couts[18][12] ;
wire \couts[18][11] ;
wire \couts[18][10] ;
wire \couts[17][63] ;
wire \couts[17][62] ;
wire \couts[17][61] ;
wire \couts[17][60] ;
wire \couts[17][59] ;
wire \couts[17][58] ;
wire \couts[17][57] ;
wire \couts[17][56] ;
wire \couts[17][55] ;
wire \couts[17][54] ;
wire \couts[17][53] ;
wire \couts[17][52] ;
wire \couts[17][51] ;
wire \couts[17][50] ;
wire \couts[17][49] ;
wire \couts[17][48] ;
wire \couts[17][47] ;
wire \couts[17][46] ;
wire \couts[17][45] ;
wire \couts[17][44] ;
wire \couts[17][43] ;
wire \couts[17][42] ;
wire \couts[17][41] ;
wire \couts[17][40] ;
wire \couts[17][39] ;
wire \couts[17][38] ;
wire \couts[17][37] ;
wire \couts[17][36] ;
wire \couts[17][35] ;
wire \couts[17][34] ;
wire \couts[17][33] ;
wire \couts[17][32] ;
wire \couts[17][31] ;
wire \couts[17][30] ;
wire \couts[17][29] ;
wire \couts[17][28] ;
wire \couts[17][27] ;
wire \couts[17][26] ;
wire \couts[17][25] ;
wire \couts[17][24] ;
wire \couts[17][23] ;
wire \couts[17][22] ;
wire \couts[17][21] ;
wire \couts[17][20] ;
wire \couts[17][19] ;
wire \couts[17][18] ;
wire \couts[17][17] ;
wire \couts[17][16] ;
wire \couts[17][15] ;
wire \couts[17][14] ;
wire \couts[17][13] ;
wire \couts[17][12] ;
wire \couts[17][11] ;
wire \couts[17][10] ;
wire \couts[17][9] ;
wire \couts[17][8] ;
wire \couts[17][7] ;
wire \couts[17][6] ;
wire \couts[17][5] ;
wire \couts[17][4] ;
wire \sums[17][63] ;
wire \sums[17][62] ;
wire \sums[17][61] ;
wire \sums[17][60] ;
wire \sums[17][59] ;
wire \sums[17][58] ;
wire \sums[17][57] ;
wire \sums[17][56] ;
wire \sums[17][55] ;
wire \sums[17][54] ;
wire \sums[17][53] ;
wire \sums[17][52] ;
wire \sums[17][51] ;
wire \sums[17][50] ;
wire \sums[17][49] ;
wire \sums[17][48] ;
wire \sums[17][47] ;
wire \sums[17][46] ;
wire \sums[17][45] ;
wire \sums[17][44] ;
wire \sums[17][43] ;
wire \sums[17][42] ;
wire \sums[17][41] ;
wire \sums[17][40] ;
wire \sums[17][39] ;
wire \sums[17][38] ;
wire \sums[17][37] ;
wire \sums[17][36] ;
wire \sums[17][35] ;
wire \sums[17][34] ;
wire \sums[17][33] ;
wire \sums[17][32] ;
wire \sums[17][31] ;
wire \sums[17][30] ;
wire \sums[17][29] ;
wire \sums[17][28] ;
wire \sums[17][27] ;
wire \sums[17][26] ;
wire \sums[17][25] ;
wire \sums[17][24] ;
wire \sums[17][23] ;
wire \sums[17][22] ;
wire \sums[17][21] ;
wire \sums[17][20] ;
wire \sums[17][19] ;
wire \sums[17][18] ;
wire \sums[17][17] ;
wire \sums[17][16] ;
wire \sums[17][15] ;
wire \sums[17][14] ;
wire \sums[17][13] ;
wire \sums[17][12] ;
wire \sums[17][11] ;
wire \sums[17][10] ;
wire \sums[17][9] ;
wire \sums[17][8] ;
wire \sums[17][7] ;
wire \sums[17][6] ;
wire \sums[17][5] ;
wire \sums[17][4] ;
wire \couts[10][62] ;
wire \couts[10][36] ;
wire \couts[10][35] ;
wire \couts[10][34] ;
wire \couts[10][33] ;
wire \couts[10][32] ;
wire \couts[10][31] ;
wire \couts[10][30] ;
wire \couts[10][29] ;
wire \couts[10][28] ;
wire \couts[10][27] ;
wire \couts[10][26] ;
wire \couts[10][25] ;
wire \couts[10][24] ;
wire \couts[10][23] ;
wire \couts[10][22] ;
wire \couts[10][21] ;
wire \couts[10][20] ;
wire \couts[10][19] ;
wire \couts[10][18] ;
wire \couts[10][17] ;
wire \couts[10][16] ;
wire \couts[10][15] ;
wire \couts[10][14] ;
wire \couts[10][13] ;
wire \couts[10][12] ;
wire \couts[10][11] ;
wire \couts[10][10] ;
wire \couts[10][9] ;
wire \couts[10][8] ;
wire \couts[10][7] ;
wire \couts[10][6] ;
wire \couts[10][5] ;
wire \couts[10][4] ;
wire \couts[10][3] ;
wire \sums[10][62] ;
wire \sums[10][35] ;
wire \sums[10][34] ;
wire \sums[10][33] ;
wire \sums[10][32] ;
wire \sums[10][31] ;
wire \sums[10][30] ;
wire \sums[10][29] ;
wire \sums[10][28] ;
wire \sums[10][27] ;
wire \sums[10][26] ;
wire \sums[10][25] ;
wire \sums[10][24] ;
wire \sums[10][23] ;
wire \sums[10][22] ;
wire \sums[10][21] ;
wire \sums[10][20] ;
wire \sums[10][19] ;
wire \sums[10][18] ;
wire \sums[10][17] ;
wire \sums[10][16] ;
wire \sums[10][15] ;
wire \sums[10][14] ;
wire \sums[10][13] ;
wire \sums[10][12] ;
wire \sums[10][11] ;
wire \sums[10][10] ;
wire \sums[10][9] ;
wire \sums[10][8] ;
wire \sums[10][7] ;
wire \sums[10][6] ;
wire \sums[10][5] ;
wire \sums[10][4] ;
wire \sums[10][3] ;
wire \couts[22][63] ;
wire \couts[22][62] ;
wire \couts[22][61] ;
wire \couts[22][60] ;
wire \couts[22][59] ;
wire \couts[22][58] ;
wire \couts[22][57] ;
wire \couts[22][56] ;
wire \couts[22][55] ;
wire \couts[22][54] ;
wire \couts[22][53] ;
wire \couts[22][52] ;
wire \couts[22][51] ;
wire \couts[22][50] ;
wire \couts[22][49] ;
wire \couts[22][48] ;
wire \couts[22][47] ;
wire \couts[22][46] ;
wire \couts[22][45] ;
wire \couts[22][44] ;
wire \couts[22][43] ;
wire \couts[22][42] ;
wire \couts[22][41] ;
wire \couts[22][40] ;
wire \couts[22][39] ;
wire \couts[22][38] ;
wire \couts[22][37] ;
wire \couts[22][36] ;
wire \couts[22][35] ;
wire \couts[22][34] ;
wire \couts[22][33] ;
wire \couts[22][32] ;
wire \couts[22][31] ;
wire \couts[22][30] ;
wire \couts[22][29] ;
wire \couts[22][28] ;
wire \couts[22][27] ;
wire \couts[22][26] ;
wire \couts[22][25] ;
wire \couts[22][24] ;
wire \couts[22][23] ;
wire \couts[22][22] ;
wire \couts[22][21] ;
wire \couts[22][20] ;
wire \couts[22][19] ;
wire \couts[22][18] ;
wire \couts[22][17] ;
wire \couts[22][16] ;
wire \couts[22][15] ;
wire \couts[22][14] ;
wire \couts[22][13] ;
wire \couts[22][12] ;
wire \couts[22][11] ;
wire \couts[22][10] ;
wire \couts[22][9] ;
wire \couts[22][8] ;
wire \couts[22][7] ;
wire \couts[22][6] ;
wire \couts[22][5] ;
wire \sums[22][63] ;
wire \sums[22][62] ;
wire \sums[22][61] ;
wire \sums[22][60] ;
wire \sums[22][59] ;
wire \sums[22][58] ;
wire \sums[22][57] ;
wire \sums[22][56] ;
wire \sums[22][55] ;
wire \sums[22][54] ;
wire \sums[22][53] ;
wire \sums[22][52] ;
wire \sums[22][51] ;
wire \sums[22][50] ;
wire \sums[22][49] ;
wire \sums[22][48] ;
wire \sums[22][47] ;
wire \sums[22][46] ;
wire \sums[22][45] ;
wire \sums[22][44] ;
wire \sums[22][43] ;
wire \sums[22][42] ;
wire \sums[22][41] ;
wire \sums[22][40] ;
wire \sums[22][39] ;
wire \sums[22][38] ;
wire \sums[22][37] ;
wire \sums[22][36] ;
wire \sums[22][35] ;
wire \sums[22][34] ;
wire \sums[22][33] ;
wire \sums[22][32] ;
wire \sums[22][31] ;
wire \sums[22][30] ;
wire \sums[22][29] ;
wire \sums[22][28] ;
wire \sums[22][27] ;
wire \sums[22][26] ;
wire \sums[22][25] ;
wire \sums[22][24] ;
wire \sums[22][23] ;
wire \sums[22][22] ;
wire \sums[22][21] ;
wire \sums[22][20] ;
wire \sums[22][19] ;
wire \sums[22][18] ;
wire \sums[22][17] ;
wire \sums[22][16] ;
wire \sums[22][15] ;
wire \sums[22][14] ;
wire \sums[22][13] ;
wire \sums[22][12] ;
wire \sums[22][11] ;
wire \sums[22][10] ;
wire \sums[22][9] ;
wire \sums[22][8] ;
wire \sums[22][7] ;
wire \sums[22][6] ;
wire \sums[22][5] ;
wire n_2_0;
wire \couts[1][37] ;
wire \couts[1][36] ;
wire \couts[1][35] ;
wire \couts[1][34] ;
wire \couts[1][33] ;
wire \couts[1][32] ;
wire \couts[1][31] ;
wire \couts[1][30] ;
wire \couts[1][29] ;
wire \couts[1][28] ;
wire \couts[1][27] ;
wire \couts[1][26] ;
wire \couts[1][25] ;
wire \couts[1][24] ;
wire \couts[1][23] ;
wire \couts[1][22] ;
wire \couts[1][21] ;
wire \couts[1][20] ;
wire \couts[1][19] ;
wire \couts[1][18] ;
wire \couts[1][17] ;
wire \couts[1][16] ;
wire \couts[1][15] ;
wire \couts[1][14] ;
wire \couts[1][13] ;
wire \couts[1][12] ;
wire \couts[1][11] ;
wire \couts[1][10] ;
wire \couts[1][9] ;
wire \couts[1][8] ;
wire \couts[1][7] ;
wire \couts[1][6] ;
wire \sums[1][61] ;
wire \sums[1][35] ;
wire \sums[1][34] ;
wire \sums[1][33] ;
wire \sums[1][32] ;
wire \sums[1][31] ;
wire \sums[1][30] ;
wire \sums[1][29] ;
wire \sums[1][28] ;
wire \sums[1][27] ;
wire \sums[1][26] ;
wire \sums[1][25] ;
wire \sums[1][24] ;
wire \sums[1][23] ;
wire \sums[1][22] ;
wire \sums[1][21] ;
wire \sums[1][20] ;
wire \sums[1][19] ;
wire \sums[1][18] ;
wire \sums[1][17] ;
wire \sums[1][16] ;
wire \sums[1][15] ;
wire \sums[1][14] ;
wire \sums[1][13] ;
wire \sums[1][12] ;
wire \sums[1][11] ;
wire \sums[1][10] ;
wire \sums[1][9] ;
wire \sums[1][8] ;
wire \sums[1][7] ;
wire \sums[1][6] ;
wire \sums[1][5] ;
wire \sums[1][4] ;
wire \couts[0][61] ;
wire \couts[0][33] ;
wire \couts[0][32] ;
wire \couts[0][31] ;
wire \couts[0][30] ;
wire \couts[0][29] ;
wire \couts[0][28] ;
wire \couts[0][27] ;
wire \couts[0][26] ;
wire \couts[0][25] ;
wire \couts[0][24] ;
wire \couts[0][23] ;
wire \couts[0][22] ;
wire \couts[0][21] ;
wire \couts[0][20] ;
wire \couts[0][19] ;
wire \couts[0][18] ;
wire \couts[0][17] ;
wire \couts[0][16] ;
wire \couts[0][15] ;
wire \couts[0][14] ;
wire \couts[0][13] ;
wire \couts[0][12] ;
wire \couts[0][11] ;
wire \couts[0][10] ;
wire \couts[0][9] ;
wire \couts[0][8] ;
wire \couts[0][7] ;
wire \couts[0][6] ;
wire \couts[0][5] ;
wire \couts[0][4] ;
wire \couts[0][3] ;
wire \couts[0][2] ;
wire \sums[0][61] ;
wire \sums[0][32] ;
wire \sums[0][31] ;
wire \sums[0][30] ;
wire \sums[0][29] ;
wire \sums[0][28] ;
wire \sums[0][27] ;
wire \sums[0][26] ;
wire \sums[0][25] ;
wire \sums[0][24] ;
wire \sums[0][23] ;
wire \sums[0][22] ;
wire \sums[0][21] ;
wire \sums[0][20] ;
wire \sums[0][19] ;
wire \sums[0][18] ;
wire \sums[0][17] ;
wire \sums[0][16] ;
wire \sums[0][15] ;
wire \sums[0][14] ;
wire \sums[0][13] ;
wire \sums[0][12] ;
wire \sums[0][11] ;
wire \sums[0][10] ;
wire \sums[0][9] ;
wire \sums[0][8] ;
wire \sums[0][7] ;
wire \sums[0][6] ;
wire \sums[0][5] ;
wire \sums[0][4] ;
wire \sums[0][3] ;
wire \sums[0][2] ;
wire \couts[25][63] ;
wire \couts[25][62] ;
wire \couts[25][61] ;
wire \couts[25][60] ;
wire \couts[25][59] ;
wire \couts[25][58] ;
wire \couts[25][57] ;
wire \couts[25][56] ;
wire \couts[25][55] ;
wire \couts[25][54] ;
wire \couts[25][53] ;
wire \couts[25][52] ;
wire \couts[25][51] ;
wire \couts[25][50] ;
wire \couts[25][49] ;
wire \couts[25][48] ;
wire \couts[25][47] ;
wire \couts[25][46] ;
wire \couts[25][45] ;
wire \couts[25][44] ;
wire \couts[25][43] ;
wire \couts[25][42] ;
wire \couts[25][41] ;
wire \couts[25][40] ;
wire \couts[25][39] ;
wire \couts[25][38] ;
wire \couts[25][37] ;
wire \couts[25][36] ;
wire \couts[25][35] ;
wire \couts[25][34] ;
wire \couts[25][33] ;
wire \couts[25][32] ;
wire \couts[25][31] ;
wire \couts[25][30] ;
wire \couts[25][29] ;
wire \couts[25][28] ;
wire \couts[25][27] ;
wire \couts[25][26] ;
wire \couts[25][25] ;
wire \couts[25][24] ;
wire \couts[25][23] ;
wire \couts[25][22] ;
wire \couts[25][21] ;
wire \couts[25][20] ;
wire \couts[25][19] ;
wire \couts[25][18] ;
wire \couts[25][17] ;
wire \couts[25][16] ;
wire \couts[25][15] ;
wire \couts[25][14] ;
wire \couts[25][13] ;
wire \couts[25][12] ;
wire \couts[25][11] ;
wire \couts[25][10] ;
wire \couts[25][9] ;
wire \couts[25][8] ;
wire \couts[25][7] ;
wire \couts[25][6] ;
wire \sums[25][63] ;
wire \sums[25][62] ;
wire \sums[25][61] ;
wire \sums[25][60] ;
wire \sums[25][59] ;
wire \sums[25][58] ;
wire \sums[25][57] ;
wire \sums[25][56] ;
wire \sums[25][55] ;
wire \sums[25][54] ;
wire \sums[25][53] ;
wire \sums[25][52] ;
wire \sums[25][51] ;
wire \sums[25][50] ;
wire \sums[25][49] ;
wire \sums[25][48] ;
wire \sums[25][47] ;
wire \sums[25][46] ;
wire \sums[25][45] ;
wire \sums[25][44] ;
wire \sums[25][43] ;
wire \sums[25][42] ;
wire \sums[25][41] ;
wire \sums[25][40] ;
wire \sums[25][39] ;
wire \sums[25][38] ;
wire \sums[25][37] ;
wire \sums[25][36] ;
wire \sums[25][35] ;
wire \sums[25][34] ;
wire \sums[25][33] ;
wire \sums[25][32] ;
wire \sums[25][31] ;
wire \sums[25][30] ;
wire \sums[25][29] ;
wire \sums[25][28] ;
wire \sums[25][27] ;
wire \sums[25][26] ;
wire \sums[25][25] ;
wire \sums[25][24] ;
wire \sums[25][23] ;
wire \sums[25][22] ;
wire \sums[25][21] ;
wire \sums[25][20] ;
wire \sums[25][19] ;
wire \sums[25][18] ;
wire \sums[25][17] ;
wire \sums[25][16] ;
wire \sums[25][15] ;
wire \sums[25][14] ;
wire \sums[25][13] ;
wire \sums[25][12] ;
wire \sums[25][11] ;
wire \sums[25][10] ;
wire \sums[25][9] ;
wire \sums[25][8] ;
wire \sums[25][7] ;
wire \sums[25][6] ;
wire \couts[7][63] ;
wire \couts[7][54] ;
wire \couts[7][53] ;
wire \couts[7][52] ;
wire \couts[7][51] ;
wire \couts[7][50] ;
wire \couts[7][49] ;
wire \couts[7][48] ;
wire \couts[7][47] ;
wire \couts[7][46] ;
wire \couts[7][45] ;
wire \couts[7][44] ;
wire \couts[7][43] ;
wire \couts[7][42] ;
wire \couts[7][41] ;
wire \couts[7][40] ;
wire \couts[7][39] ;
wire \couts[7][38] ;
wire \couts[7][37] ;
wire \couts[7][36] ;
wire \couts[7][35] ;
wire \couts[7][34] ;
wire \couts[7][33] ;
wire \couts[7][32] ;
wire \couts[7][31] ;
wire \couts[7][30] ;
wire \couts[7][29] ;
wire \couts[7][28] ;
wire \couts[7][27] ;
wire \couts[7][26] ;
wire \couts[7][25] ;
wire \couts[7][24] ;
wire \couts[7][23] ;
wire \sums[7][63] ;
wire \sums[7][53] ;
wire \sums[7][52] ;
wire \sums[7][51] ;
wire \sums[7][50] ;
wire \sums[7][49] ;
wire \sums[7][48] ;
wire \sums[7][47] ;
wire \sums[7][46] ;
wire \sums[7][45] ;
wire \sums[7][44] ;
wire \sums[7][43] ;
wire \sums[7][42] ;
wire \sums[7][41] ;
wire \sums[7][40] ;
wire \sums[7][39] ;
wire \sums[7][38] ;
wire \sums[7][37] ;
wire \sums[7][36] ;
wire \sums[7][35] ;
wire \sums[7][34] ;
wire \sums[7][33] ;
wire \sums[7][32] ;
wire \sums[7][31] ;
wire \sums[7][30] ;
wire \sums[7][29] ;
wire \sums[7][28] ;
wire \sums[7][27] ;
wire \sums[7][26] ;
wire \sums[7][25] ;
wire \sums[7][24] ;
wire \sums[7][23] ;
wire \sums[7][22] ;
wire \sums[20][59] ;
wire \sums[20][58] ;
wire \sums[20][57] ;
wire \sums[20][56] ;
wire \sums[20][55] ;
wire \sums[20][54] ;
wire \sums[20][53] ;
wire \sums[20][52] ;
wire \sums[20][51] ;
wire \sums[20][50] ;
wire \sums[20][49] ;
wire \sums[20][48] ;
wire \sums[20][47] ;
wire \sums[20][46] ;
wire \sums[20][45] ;
wire \sums[20][44] ;
wire \sums[20][43] ;
wire \sums[20][42] ;
wire \sums[20][41] ;
wire \sums[20][40] ;
wire \sums[20][39] ;
wire \sums[20][38] ;
wire \sums[20][37] ;
wire \sums[20][36] ;
wire \sums[20][35] ;
wire \sums[20][34] ;
wire \sums[20][33] ;
wire \sums[20][32] ;
wire \sums[20][31] ;
wire \sums[20][30] ;
wire \sums[20][29] ;
wire \sums[20][28] ;
wire \sums[20][27] ;
wire \sums[20][26] ;
wire \sums[20][25] ;
wire \sums[20][24] ;
wire \sums[20][23] ;
wire \sums[20][22] ;
wire \sums[20][21] ;
wire \couts[14][63] ;
wire \couts[14][54] ;
wire \couts[14][53] ;
wire \couts[14][52] ;
wire \couts[14][51] ;
wire \couts[14][50] ;
wire \couts[14][49] ;
wire \couts[14][48] ;
wire \couts[14][47] ;
wire \couts[14][46] ;
wire \couts[14][45] ;
wire \couts[14][44] ;
wire \couts[14][43] ;
wire \couts[14][42] ;
wire \couts[14][41] ;
wire \couts[14][40] ;
wire \couts[14][39] ;
wire \couts[14][38] ;
wire \couts[14][37] ;
wire \couts[14][36] ;
wire \couts[14][35] ;
wire \couts[14][34] ;
wire \couts[14][33] ;
wire \couts[14][32] ;
wire \couts[14][31] ;
wire \couts[14][30] ;
wire \couts[14][29] ;
wire \couts[14][28] ;
wire \couts[14][27] ;
wire \couts[14][26] ;
wire \couts[14][25] ;
wire \couts[14][24] ;
wire \couts[14][23] ;
wire \sums[14][63] ;
wire \sums[14][53] ;
wire \sums[14][52] ;
wire \sums[14][51] ;
wire \sums[14][50] ;
wire \sums[14][49] ;
wire \sums[14][48] ;
wire \sums[14][47] ;
wire \sums[14][46] ;
wire \sums[14][45] ;
wire \sums[14][44] ;
wire \sums[14][43] ;
wire \sums[14][42] ;
wire \sums[14][41] ;
wire \sums[14][40] ;
wire \sums[14][39] ;
wire \sums[14][38] ;
wire \sums[14][37] ;
wire \sums[14][36] ;
wire \sums[14][35] ;
wire \sums[14][34] ;
wire \sums[14][33] ;
wire \sums[14][32] ;
wire \sums[14][31] ;
wire \sums[14][30] ;
wire \sums[14][29] ;
wire \sums[14][28] ;
wire \sums[14][27] ;
wire \sums[14][26] ;
wire \sums[14][25] ;
wire \sums[14][24] ;
wire \sums[14][23] ;
wire \sums[14][22] ;
wire \sums[14][21] ;
wire \sums[14][20] ;
wire \couts[19][63] ;
wire \couts[19][54] ;
wire \couts[19][53] ;
wire \couts[19][52] ;
wire \couts[19][51] ;
wire \couts[19][50] ;
wire \couts[19][49] ;
wire \couts[19][48] ;
wire \couts[19][47] ;
wire \couts[19][46] ;
wire \couts[19][45] ;
wire \couts[19][44] ;
wire \couts[19][43] ;
wire \couts[19][42] ;
wire \couts[19][41] ;
wire \couts[19][40] ;
wire \couts[19][39] ;
wire \couts[19][38] ;
wire \couts[19][37] ;
wire \couts[19][36] ;
wire \couts[19][35] ;
wire \couts[19][34] ;
wire \couts[19][33] ;
wire \couts[19][32] ;
wire \couts[19][31] ;
wire \couts[19][30] ;
wire \couts[19][29] ;
wire \couts[19][28] ;
wire \couts[19][27] ;
wire \couts[19][26] ;
wire \couts[19][25] ;
wire \couts[19][24] ;
wire \couts[19][23] ;
wire \couts[19][22] ;
wire \couts[19][21] ;
wire \couts[19][20] ;
wire \couts[19][19] ;
wire \couts[19][18] ;
wire \couts[19][17] ;
wire \sums[19][63] ;
wire \sums[19][53] ;
wire \sums[19][52] ;
wire \sums[19][51] ;
wire \sums[19][50] ;
wire \sums[19][49] ;
wire \sums[19][48] ;
wire \sums[19][47] ;
wire \sums[19][46] ;
wire \sums[19][45] ;
wire \sums[19][44] ;
wire \sums[19][43] ;
wire \sums[19][42] ;
wire \sums[19][41] ;
wire \sums[19][40] ;
wire \sums[19][39] ;
wire \sums[19][38] ;
wire \sums[19][37] ;
wire \sums[19][36] ;
wire \sums[19][35] ;
wire \sums[19][34] ;
wire \sums[19][33] ;
wire \sums[19][32] ;
wire \sums[19][31] ;
wire \sums[19][30] ;
wire \sums[19][29] ;
wire \sums[19][28] ;
wire \sums[19][27] ;
wire \sums[19][26] ;
wire \sums[19][25] ;
wire \sums[19][24] ;
wire \sums[19][23] ;
wire \sums[19][22] ;
wire \sums[19][21] ;
wire \sums[19][20] ;
wire \sums[19][19] ;
wire \sums[19][18] ;
wire \sums[19][17] ;
wire \sums[19][16] ;
wire \couts[23][63] ;
wire \couts[23][62] ;
wire \couts[23][61] ;
wire \couts[23][60] ;
wire \couts[23][59] ;
wire \couts[23][58] ;
wire \couts[23][57] ;
wire \couts[23][56] ;
wire \couts[23][55] ;
wire \couts[23][54] ;
wire \couts[23][53] ;
wire \couts[23][52] ;
wire \couts[23][51] ;
wire \couts[23][50] ;
wire \couts[23][49] ;
wire \couts[23][48] ;
wire \couts[23][47] ;
wire \couts[23][46] ;
wire \couts[23][45] ;
wire \couts[23][44] ;
wire \couts[23][43] ;
wire \couts[23][42] ;
wire \couts[23][41] ;
wire \couts[23][40] ;
wire \couts[23][39] ;
wire \couts[23][38] ;
wire \couts[23][37] ;
wire \couts[23][36] ;
wire \couts[23][35] ;
wire \couts[23][34] ;
wire \couts[23][33] ;
wire \couts[23][32] ;
wire \couts[23][31] ;
wire \couts[23][30] ;
wire \couts[23][29] ;
wire \couts[23][28] ;
wire \couts[23][27] ;
wire \couts[23][26] ;
wire \couts[23][25] ;
wire \couts[23][24] ;
wire \couts[23][23] ;
wire \couts[23][22] ;
wire \couts[23][21] ;
wire \couts[23][20] ;
wire \couts[23][19] ;
wire \couts[23][18] ;
wire \couts[23][17] ;
wire \couts[23][16] ;
wire \couts[23][15] ;
wire \sums[23][63] ;
wire \sums[23][62] ;
wire \sums[23][61] ;
wire \sums[23][60] ;
wire \sums[23][59] ;
wire \sums[23][58] ;
wire \sums[23][57] ;
wire \sums[23][56] ;
wire \sums[23][55] ;
wire \sums[23][54] ;
wire \sums[23][53] ;
wire \sums[23][52] ;
wire \sums[23][51] ;
wire \sums[23][50] ;
wire \sums[23][49] ;
wire \sums[23][48] ;
wire \sums[23][47] ;
wire \sums[23][46] ;
wire \sums[23][45] ;
wire \sums[23][44] ;
wire \sums[23][43] ;
wire \sums[23][42] ;
wire \sums[23][41] ;
wire \sums[23][40] ;
wire \sums[23][39] ;
wire \sums[23][38] ;
wire \sums[23][37] ;
wire \sums[23][36] ;
wire \sums[23][35] ;
wire \sums[23][34] ;
wire \sums[23][33] ;
wire \sums[23][32] ;
wire \sums[23][31] ;
wire \sums[23][30] ;
wire \sums[23][29] ;
wire \sums[23][28] ;
wire \sums[23][27] ;
wire \sums[23][26] ;
wire \sums[23][25] ;
wire \sums[23][24] ;
wire \sums[23][23] ;
wire \sums[23][22] ;
wire \sums[23][21] ;
wire \sums[23][20] ;
wire \sums[23][19] ;
wire \sums[23][18] ;
wire \sums[23][17] ;
wire \sums[23][16] ;
wire \sums[23][15] ;
wire \sums[23][14] ;
wire \couts[6][63] ;
wire \couts[6][51] ;
wire \couts[6][50] ;
wire \couts[6][49] ;
wire \couts[6][48] ;
wire \couts[6][47] ;
wire \couts[6][46] ;
wire \couts[6][45] ;
wire \couts[6][44] ;
wire \couts[6][43] ;
wire \couts[6][42] ;
wire \couts[6][41] ;
wire \couts[6][40] ;
wire \couts[6][39] ;
wire \couts[6][38] ;
wire \couts[6][37] ;
wire \couts[6][36] ;
wire \couts[6][35] ;
wire \couts[6][34] ;
wire \couts[6][33] ;
wire \couts[6][32] ;
wire \couts[6][31] ;
wire \couts[6][30] ;
wire \couts[6][29] ;
wire \couts[6][28] ;
wire \couts[6][27] ;
wire \couts[6][26] ;
wire \couts[6][25] ;
wire \couts[6][24] ;
wire \couts[6][23] ;
wire \couts[6][22] ;
wire \couts[6][21] ;
wire \couts[6][20] ;
wire \sums[6][63] ;
wire \sums[6][50] ;
wire \sums[6][49] ;
wire \sums[6][48] ;
wire \sums[6][47] ;
wire \sums[6][46] ;
wire \sums[6][45] ;
wire \sums[6][44] ;
wire \sums[6][43] ;
wire \sums[6][42] ;
wire \sums[6][41] ;
wire \sums[6][40] ;
wire \sums[6][39] ;
wire \sums[6][38] ;
wire \sums[6][37] ;
wire \sums[6][36] ;
wire \sums[6][35] ;
wire \sums[6][34] ;
wire \sums[6][33] ;
wire \sums[6][32] ;
wire \sums[6][31] ;
wire \sums[6][30] ;
wire \sums[6][29] ;
wire \sums[6][28] ;
wire \sums[6][27] ;
wire \sums[6][26] ;
wire \sums[6][25] ;
wire \sums[6][24] ;
wire \sums[6][23] ;
wire \sums[6][22] ;
wire \sums[6][21] ;
wire \sums[6][20] ;
wire \sums[6][19] ;
wire \couts[8][63] ;
wire \couts[8][57] ;
wire \couts[8][56] ;
wire \couts[8][55] ;
wire \couts[8][54] ;
wire \couts[8][53] ;
wire \couts[8][52] ;
wire \couts[8][51] ;
wire \couts[8][50] ;
wire \couts[8][49] ;
wire \couts[8][48] ;
wire \couts[8][47] ;
wire \couts[8][46] ;
wire \couts[8][45] ;
wire \couts[8][44] ;
wire \couts[8][43] ;
wire \couts[8][42] ;
wire \couts[8][41] ;
wire \couts[8][40] ;
wire \couts[8][39] ;
wire \couts[8][38] ;
wire \couts[8][37] ;
wire \couts[8][36] ;
wire \couts[8][35] ;
wire \couts[8][34] ;
wire \couts[8][33] ;
wire \couts[8][32] ;
wire \couts[8][31] ;
wire \couts[8][30] ;
wire \couts[8][29] ;
wire \couts[8][28] ;
wire \couts[8][27] ;
wire \couts[8][26] ;
wire \sums[8][63] ;
wire \sums[8][56] ;
wire \sums[8][55] ;
wire \sums[8][54] ;
wire \sums[8][53] ;
wire \sums[8][52] ;
wire \sums[8][51] ;
wire \sums[8][50] ;
wire \sums[8][49] ;
wire \sums[8][48] ;
wire \sums[8][47] ;
wire \sums[8][46] ;
wire \sums[8][45] ;
wire \sums[8][44] ;
wire \sums[8][43] ;
wire \sums[8][42] ;
wire \sums[8][41] ;
wire \sums[8][40] ;
wire \sums[8][39] ;
wire \sums[8][38] ;
wire \sums[8][37] ;
wire \sums[8][36] ;
wire \sums[8][35] ;
wire \sums[8][34] ;
wire \sums[8][33] ;
wire \sums[8][32] ;
wire \sums[8][31] ;
wire \sums[8][30] ;
wire \sums[8][29] ;
wire \sums[8][28] ;
wire \sums[8][27] ;
wire \sums[8][26] ;
wire \sums[8][25] ;
wire \couts[15][63] ;
wire \couts[15][58] ;
wire \couts[15][57] ;
wire \couts[15][56] ;
wire \couts[15][55] ;
wire \couts[15][54] ;
wire \couts[15][53] ;
wire \couts[15][52] ;
wire \couts[15][51] ;
wire \couts[15][50] ;
wire \couts[15][49] ;
wire \couts[15][48] ;
wire \couts[15][47] ;
wire \couts[15][46] ;
wire \couts[15][45] ;
wire \couts[15][44] ;
wire \couts[15][43] ;
wire \couts[15][42] ;
wire \couts[15][41] ;
wire \couts[15][40] ;
wire \couts[15][39] ;
wire \couts[15][38] ;
wire \couts[15][37] ;
wire \couts[15][36] ;
wire \couts[15][35] ;
wire \couts[15][34] ;
wire \couts[15][33] ;
wire \couts[15][32] ;
wire \couts[15][31] ;
wire \couts[15][30] ;
wire \couts[15][29] ;
wire \couts[15][28] ;
wire \couts[15][27] ;
wire \couts[15][26] ;
wire \couts[15][25] ;
wire \sums[15][63] ;
wire \sums[15][57] ;
wire \sums[15][56] ;
wire \sums[15][55] ;
wire \sums[15][54] ;
wire \sums[15][53] ;
wire \sums[15][52] ;
wire \sums[15][51] ;
wire \sums[15][50] ;
wire \sums[15][49] ;
wire \sums[15][48] ;
wire \sums[15][47] ;
wire \sums[15][46] ;
wire \sums[15][45] ;
wire \sums[15][44] ;
wire \sums[15][43] ;
wire \sums[15][42] ;
wire \sums[15][41] ;
wire \sums[15][40] ;
wire \sums[15][39] ;
wire \sums[15][38] ;
wire \sums[15][37] ;
wire \sums[15][36] ;
wire \sums[15][35] ;
wire \sums[15][34] ;
wire \sums[15][33] ;
wire \sums[15][32] ;
wire \sums[15][31] ;
wire \sums[15][30] ;
wire \sums[15][29] ;
wire \sums[15][28] ;
wire \sums[15][27] ;
wire \sums[15][26] ;
wire \sums[15][25] ;
wire \sums[15][24] ;
wire \couts[20][63] ;
wire \couts[20][59] ;
wire \couts[20][58] ;
wire \couts[20][57] ;
wire \couts[20][56] ;
wire \couts[20][55] ;
wire \couts[20][54] ;
wire \couts[20][53] ;
wire \couts[20][52] ;
wire \couts[20][51] ;
wire \couts[20][50] ;
wire \couts[20][49] ;
wire \couts[20][48] ;
wire \couts[20][47] ;
wire \couts[20][46] ;
wire \couts[20][45] ;
wire \couts[20][44] ;
wire \couts[20][43] ;
wire \couts[20][42] ;
wire \couts[20][41] ;
wire \couts[20][40] ;
wire \couts[20][39] ;
wire \couts[20][38] ;
wire \couts[20][37] ;
wire \couts[20][36] ;
wire \couts[20][35] ;
wire \couts[20][34] ;
wire \couts[20][33] ;
wire \couts[20][32] ;
wire \couts[20][31] ;
wire \couts[20][30] ;
wire \couts[20][29] ;
wire \couts[20][28] ;
wire \couts[20][27] ;
wire \couts[20][26] ;
wire \couts[20][25] ;
wire \couts[20][24] ;
wire \couts[9][63] ;
wire \couts[9][62] ;
wire \couts[9][61] ;
wire \couts[9][60] ;
wire \couts[9][59] ;
wire \couts[9][58] ;
wire \couts[9][57] ;
wire \couts[9][56] ;
wire \couts[9][55] ;
wire \couts[9][54] ;
wire \couts[9][53] ;
wire \couts[9][52] ;
wire \couts[9][51] ;
wire \couts[9][50] ;
wire \couts[9][49] ;
wire \couts[9][48] ;
wire \couts[9][47] ;
wire \couts[9][46] ;
wire \couts[9][45] ;
wire \couts[9][44] ;
wire \couts[9][43] ;
wire \couts[9][42] ;
wire \couts[9][41] ;
wire \couts[9][40] ;
wire \couts[9][39] ;
wire \couts[9][38] ;
wire \couts[9][37] ;
wire \couts[9][36] ;
wire \couts[9][35] ;
wire \couts[9][34] ;
wire \couts[9][33] ;
wire \couts[9][32] ;
wire \couts[9][31] ;
wire \couts[9][30] ;
wire \couts[9][29] ;
wire \sums[9][63] ;
wire \sums[9][62] ;
wire \sums[9][61] ;
wire \sums[9][60] ;
wire \sums[9][59] ;
wire \sums[9][58] ;
wire \sums[9][57] ;
wire \sums[9][56] ;
wire \sums[9][55] ;
wire \sums[9][54] ;
wire \sums[9][53] ;
wire \sums[9][52] ;
wire \sums[9][51] ;
wire \sums[9][50] ;
wire \sums[9][49] ;
wire \sums[9][48] ;
wire \sums[9][47] ;
wire \sums[9][46] ;
wire \sums[9][45] ;
wire \sums[9][44] ;
wire \sums[9][43] ;
wire \sums[9][42] ;
wire \sums[9][41] ;
wire \sums[9][40] ;
wire \sums[9][39] ;
wire \sums[9][38] ;
wire \sums[9][37] ;
wire \sums[9][36] ;
wire \sums[9][35] ;
wire \sums[9][34] ;
wire \sums[9][33] ;
wire \sums[9][32] ;
wire \sums[9][31] ;
wire \sums[9][30] ;
wire \sums[9][29] ;
wire \sums[9][28] ;
wire \couts[16][63] ;
wire \couts[16][62] ;
wire \couts[16][61] ;
wire \couts[16][60] ;
wire \couts[16][59] ;
wire \couts[16][58] ;
wire \couts[16][57] ;
wire \couts[16][56] ;
wire \couts[16][55] ;
wire \couts[16][54] ;
wire \couts[16][53] ;
wire \couts[16][52] ;
wire \couts[16][51] ;
wire \couts[16][50] ;
wire \couts[16][49] ;
wire \couts[16][48] ;
wire \couts[16][47] ;
wire \couts[16][46] ;
wire \couts[16][45] ;
wire \couts[16][44] ;
wire \couts[16][43] ;
wire \couts[16][42] ;
wire \couts[16][41] ;
wire \couts[16][40] ;
wire \couts[16][39] ;
wire \couts[16][38] ;
wire \couts[16][37] ;
wire \couts[16][36] ;
wire \couts[16][35] ;
wire \couts[16][34] ;
wire \couts[16][33] ;
wire \couts[16][32] ;
wire \couts[16][31] ;
wire \couts[16][30] ;
wire \sums[16][63] ;
wire \sums[16][62] ;
wire \sums[16][61] ;
wire \sums[16][60] ;
wire \sums[16][59] ;
wire \sums[16][58] ;
wire \sums[16][57] ;
wire \sums[16][56] ;
wire \sums[16][55] ;
wire \sums[16][54] ;
wire \sums[16][53] ;
wire \sums[16][52] ;
wire \sums[16][51] ;
wire \sums[16][50] ;
wire \sums[16][49] ;
wire \sums[16][48] ;
wire \sums[16][47] ;
wire \sums[16][46] ;
wire \sums[16][45] ;
wire \sums[16][44] ;
wire \sums[16][43] ;
wire \sums[16][42] ;
wire \sums[16][41] ;
wire \sums[16][40] ;
wire \sums[16][39] ;
wire \sums[16][38] ;
wire \sums[16][37] ;
wire \sums[16][36] ;
wire \sums[16][35] ;
wire \sums[16][34] ;
wire \sums[16][33] ;
wire \sums[16][32] ;
wire \sums[16][31] ;
wire \sums[16][30] ;
wire \sums[16][29] ;
wire \couts[21][63] ;
wire \couts[21][62] ;
wire \couts[21][61] ;
wire \couts[21][60] ;
wire \couts[21][59] ;
wire \couts[21][58] ;
wire \couts[21][57] ;
wire \couts[21][56] ;
wire \couts[21][55] ;
wire \couts[21][54] ;
wire \couts[21][53] ;
wire \couts[21][52] ;
wire \couts[21][51] ;
wire \couts[21][50] ;
wire \couts[21][49] ;
wire \couts[21][48] ;
wire \couts[21][47] ;
wire \couts[21][46] ;
wire \couts[21][45] ;
wire \couts[21][44] ;
wire \couts[21][43] ;
wire \couts[21][42] ;
wire \couts[21][41] ;
wire \couts[21][40] ;
wire \couts[21][39] ;
wire \couts[21][38] ;
wire \couts[21][37] ;
wire \couts[21][36] ;
wire \couts[21][35] ;
wire \couts[21][34] ;
wire \couts[21][33] ;
wire \couts[21][32] ;
wire \couts[21][31] ;
wire \sums[21][63] ;
wire \sums[21][62] ;
wire \sums[21][61] ;
wire \sums[21][60] ;
wire \sums[21][59] ;
wire \sums[21][58] ;
wire \sums[21][57] ;
wire \sums[21][56] ;
wire \sums[21][55] ;
wire \sums[21][54] ;
wire \sums[21][53] ;
wire \sums[21][52] ;
wire \sums[21][51] ;
wire \sums[21][50] ;
wire \sums[21][49] ;
wire \sums[21][48] ;
wire \sums[21][47] ;
wire \sums[21][46] ;
wire \sums[21][45] ;
wire \sums[21][44] ;
wire \sums[21][43] ;
wire \sums[21][42] ;
wire \sums[21][41] ;
wire \sums[21][40] ;
wire \sums[21][39] ;
wire \sums[21][38] ;
wire \sums[21][37] ;
wire \sums[21][36] ;
wire \sums[21][35] ;
wire \sums[21][34] ;
wire \sums[21][33] ;
wire \sums[21][32] ;
wire \sums[21][31] ;
wire \sums[21][30] ;
wire \couts[24][63] ;
wire \couts[24][62] ;
wire \couts[24][61] ;
wire \couts[24][60] ;
wire \couts[24][59] ;
wire \couts[24][58] ;
wire \couts[24][57] ;
wire \couts[24][56] ;
wire \couts[24][55] ;
wire \couts[24][54] ;
wire \couts[24][53] ;
wire \couts[24][52] ;
wire \couts[24][51] ;
wire \couts[24][50] ;
wire \couts[24][49] ;
wire \couts[24][48] ;
wire \couts[24][47] ;
wire \couts[24][46] ;
wire \couts[24][45] ;
wire \couts[24][44] ;
wire \couts[24][43] ;
wire \couts[24][42] ;
wire \couts[24][41] ;
wire \couts[24][40] ;
wire \couts[24][39] ;
wire \couts[24][38] ;
wire \couts[24][37] ;
wire \couts[24][36] ;
wire \couts[24][35] ;
wire \couts[24][34] ;
wire \couts[24][33] ;
wire \couts[24][32] ;
wire \couts[24][31] ;
wire \couts[24][30] ;
wire \couts[24][29] ;
wire \couts[24][28] ;
wire \couts[24][27] ;
wire \couts[24][26] ;
wire \couts[24][25] ;
wire \sums[24][63] ;
wire \sums[24][62] ;
wire \sums[24][61] ;
wire \sums[24][60] ;
wire \sums[24][59] ;
wire \sums[24][58] ;
wire \sums[24][57] ;
wire \sums[24][56] ;
wire \sums[24][55] ;
wire \sums[24][54] ;
wire \sums[24][53] ;
wire \sums[24][52] ;
wire \sums[24][51] ;
wire \sums[24][50] ;
wire \sums[24][49] ;
wire \sums[24][48] ;
wire \sums[24][47] ;
wire \sums[24][46] ;
wire \sums[24][45] ;
wire \sums[24][44] ;
wire \sums[24][43] ;
wire \sums[24][42] ;
wire \sums[24][41] ;
wire \sums[24][40] ;
wire \sums[24][39] ;
wire \sums[24][38] ;
wire \sums[24][37] ;
wire \sums[24][36] ;
wire \sums[24][35] ;
wire \sums[24][34] ;
wire \sums[24][33] ;
wire \sums[24][32] ;
wire \sums[24][31] ;
wire \sums[24][30] ;
wire \sums[24][29] ;
wire \sums[24][28] ;
wire \sums[24][27] ;
wire \sums[24][26] ;
wire \sums[24][25] ;
wire \sums[24][24] ;
wire \couts[26][63] ;
wire \couts[26][62] ;
wire \couts[26][61] ;
wire \couts[26][60] ;
wire \couts[26][59] ;
wire \couts[26][58] ;
wire \couts[26][57] ;
wire \couts[26][56] ;
wire \couts[26][55] ;
wire \couts[26][54] ;
wire \couts[26][53] ;
wire \couts[26][52] ;
wire \couts[26][51] ;
wire \couts[26][50] ;
wire \couts[26][49] ;
wire \couts[26][48] ;
wire \couts[26][47] ;
wire \couts[26][46] ;
wire \couts[26][45] ;
wire \couts[26][44] ;
wire \couts[26][43] ;
wire \couts[26][42] ;
wire \couts[26][41] ;
wire \couts[26][40] ;
wire \couts[26][39] ;
wire \couts[26][38] ;
wire \couts[26][37] ;
wire \couts[26][36] ;
wire \couts[26][35] ;
wire \couts[26][34] ;
wire \couts[26][33] ;
wire \couts[26][32] ;
wire \couts[26][31] ;
wire \couts[26][30] ;
wire \couts[26][29] ;
wire \couts[26][28] ;
wire \couts[26][27] ;
wire \couts[26][26] ;
wire \couts[26][25] ;
wire \couts[26][24] ;
wire \couts[26][23] ;
wire \couts[26][22] ;
wire \sums[26][63] ;
wire \sums[26][62] ;
wire \sums[26][61] ;
wire \sums[26][60] ;
wire \sums[26][59] ;
wire \sums[26][58] ;
wire \sums[26][57] ;
wire \sums[26][56] ;
wire \sums[26][55] ;
wire \sums[26][54] ;
wire \sums[26][53] ;
wire \sums[26][52] ;
wire \sums[26][51] ;
wire \sums[26][50] ;
wire \sums[26][49] ;
wire \sums[26][48] ;
wire \sums[26][47] ;
wire \sums[26][46] ;
wire \sums[26][45] ;
wire \sums[26][44] ;
wire \sums[26][43] ;
wire \sums[26][42] ;
wire \sums[26][41] ;
wire \sums[26][40] ;
wire \sums[26][39] ;
wire \sums[26][38] ;
wire \sums[26][37] ;
wire \sums[26][36] ;
wire \sums[26][35] ;
wire \sums[26][34] ;
wire \sums[26][33] ;
wire \sums[26][32] ;
wire \sums[26][31] ;
wire \sums[26][30] ;
wire \sums[26][29] ;
wire \sums[26][28] ;
wire \sums[26][27] ;
wire \sums[26][26] ;
wire \sums[26][25] ;
wire \sums[26][24] ;
wire \sums[26][23] ;
wire \sums[26][22] ;
wire \sums[26][21] ;
wire \couts[27][63] ;
wire \couts[27][62] ;
wire \couts[27][61] ;
wire \couts[27][60] ;
wire \couts[27][59] ;
wire \couts[27][58] ;
wire \couts[27][57] ;
wire \couts[27][56] ;
wire \couts[27][55] ;
wire \couts[27][54] ;
wire \couts[27][53] ;
wire \couts[27][52] ;
wire \couts[27][51] ;
wire \couts[27][50] ;
wire \couts[27][49] ;
wire \couts[27][48] ;
wire \couts[27][47] ;
wire \couts[27][46] ;
wire \couts[27][45] ;
wire \couts[27][44] ;
wire \couts[27][43] ;
wire \couts[27][42] ;
wire \couts[27][41] ;
wire \couts[27][40] ;
wire \couts[27][39] ;
wire \couts[27][38] ;
wire \couts[27][37] ;
wire \couts[27][36] ;
wire \couts[27][35] ;
wire \couts[27][34] ;
wire \couts[27][33] ;
wire \couts[27][32] ;
wire \couts[27][31] ;
wire \couts[27][30] ;
wire \couts[27][29] ;
wire \couts[27][28] ;
wire \couts[27][27] ;
wire \couts[27][26] ;
wire \couts[27][25] ;
wire \couts[27][24] ;
wire \couts[27][23] ;
wire \couts[27][22] ;
wire \couts[27][21] ;
wire \couts[27][20] ;
wire \couts[27][19] ;
wire \couts[27][18] ;
wire \couts[27][17] ;
wire \couts[27][16] ;
wire \couts[27][15] ;
wire \couts[27][14] ;
wire \couts[27][13] ;
wire \couts[27][12] ;
wire \couts[27][11] ;
wire \couts[27][10] ;
wire \couts[27][9] ;
wire \couts[27][8] ;
wire \couts[27][7] ;
wire \sums[27][63] ;
wire \sums[27][62] ;
wire \sums[27][61] ;
wire \sums[27][60] ;
wire \sums[27][59] ;
wire \sums[27][58] ;
wire \sums[27][57] ;
wire \sums[27][56] ;
wire \sums[27][55] ;
wire \sums[27][54] ;
wire \sums[27][53] ;
wire \sums[27][52] ;
wire \sums[27][51] ;
wire \sums[27][50] ;
wire \sums[27][49] ;
wire \sums[27][48] ;
wire \sums[27][47] ;
wire \sums[27][46] ;
wire \sums[27][45] ;
wire \sums[27][44] ;
wire \sums[27][43] ;
wire \sums[27][42] ;
wire \sums[27][41] ;
wire \sums[27][40] ;
wire \sums[27][39] ;
wire \sums[27][38] ;
wire \sums[27][37] ;
wire \sums[27][36] ;
wire \sums[27][35] ;
wire \sums[27][34] ;
wire \sums[27][33] ;
wire \sums[27][32] ;
wire \sums[27][31] ;
wire \sums[27][30] ;
wire \sums[27][29] ;
wire \sums[27][28] ;
wire \sums[27][27] ;
wire \sums[27][26] ;
wire \sums[27][25] ;
wire \sums[27][24] ;
wire \sums[27][23] ;
wire \sums[27][22] ;
wire \sums[27][21] ;
wire \sums[27][20] ;
wire \sums[27][19] ;
wire \sums[27][18] ;
wire \sums[27][17] ;
wire \sums[27][16] ;
wire \sums[27][15] ;
wire \sums[27][14] ;
wire \sums[27][13] ;
wire \sums[27][12] ;
wire \sums[27][11] ;
wire \sums[27][10] ;
wire \sums[27][9] ;
wire \sums[27][8] ;
wire \sums[27][7] ;
wire \couts[28][63] ;
wire \couts[28][62] ;
wire \couts[28][61] ;
wire \couts[28][60] ;
wire \couts[28][59] ;
wire \couts[28][58] ;
wire \couts[28][57] ;
wire \couts[28][56] ;
wire \couts[28][55] ;
wire \couts[28][54] ;
wire \couts[28][53] ;
wire \couts[28][52] ;
wire \couts[28][51] ;
wire \couts[28][50] ;
wire \couts[28][49] ;
wire \couts[28][48] ;
wire \couts[28][47] ;
wire \couts[28][46] ;
wire \couts[28][45] ;
wire \couts[28][44] ;
wire \couts[28][43] ;
wire \couts[28][42] ;
wire \couts[28][41] ;
wire \couts[28][40] ;
wire \couts[28][39] ;
wire \couts[28][38] ;
wire \couts[28][37] ;
wire \couts[28][36] ;
wire \couts[28][35] ;
wire \couts[28][34] ;
wire \couts[28][33] ;
wire \couts[28][32] ;
wire \couts[28][31] ;
wire \couts[28][30] ;
wire \couts[28][29] ;
wire \couts[28][28] ;
wire \couts[28][27] ;
wire \couts[28][26] ;
wire \couts[28][25] ;
wire \couts[28][24] ;
wire \couts[28][23] ;
wire \couts[28][22] ;
wire \couts[28][21] ;
wire \couts[28][20] ;
wire \couts[28][19] ;
wire \couts[28][18] ;
wire \couts[28][17] ;
wire \couts[28][16] ;
wire \couts[28][15] ;
wire \couts[28][14] ;
wire \couts[28][13] ;
wire \couts[28][12] ;
wire \couts[28][11] ;
wire \couts[28][10] ;
wire \couts[28][9] ;
wire \couts[28][8] ;
wire \sums[28][63] ;
wire \sums[28][62] ;
wire \sums[28][61] ;
wire \sums[28][60] ;
wire \sums[28][59] ;
wire \sums[28][58] ;
wire \sums[28][57] ;
wire \sums[28][56] ;
wire \sums[28][55] ;
wire \sums[28][54] ;
wire \sums[28][53] ;
wire \sums[28][52] ;
wire \sums[28][51] ;
wire \sums[28][50] ;
wire \sums[28][49] ;
wire \sums[28][48] ;
wire \sums[28][47] ;
wire \sums[28][46] ;
wire \sums[28][45] ;
wire \sums[28][44] ;
wire \sums[28][43] ;
wire \sums[28][42] ;
wire \sums[28][41] ;
wire \sums[28][40] ;
wire \sums[28][39] ;
wire \sums[28][38] ;
wire \sums[28][37] ;
wire \sums[28][36] ;
wire \sums[28][35] ;
wire \sums[28][34] ;
wire \sums[28][33] ;
wire \sums[28][32] ;
wire \sums[28][31] ;
wire \sums[28][30] ;
wire \sums[28][29] ;
wire \sums[28][28] ;
wire \sums[28][27] ;
wire \sums[28][26] ;
wire \sums[28][25] ;
wire \sums[28][24] ;
wire \sums[28][23] ;
wire \sums[28][22] ;
wire \sums[28][21] ;
wire \sums[28][20] ;
wire \sums[28][19] ;
wire \sums[28][18] ;
wire \sums[28][17] ;
wire \sums[28][16] ;
wire \sums[28][15] ;
wire \sums[28][14] ;
wire \sums[28][13] ;
wire \sums[28][12] ;
wire \sums[28][11] ;
wire \sums[28][10] ;
wire \sums[28][9] ;
wire \sums[28][8] ;
wire \couts[29][63] ;
wire \couts[29][62] ;
wire \couts[29][61] ;
wire \couts[29][60] ;
wire \couts[29][59] ;
wire \couts[29][58] ;
wire \couts[29][57] ;
wire \couts[29][56] ;
wire \couts[29][55] ;
wire \couts[29][54] ;
wire \couts[29][53] ;
wire \couts[29][52] ;
wire \couts[29][51] ;
wire \couts[29][50] ;
wire \couts[29][49] ;
wire \couts[29][48] ;
wire \couts[29][47] ;
wire \couts[29][46] ;
wire \couts[29][45] ;
wire \couts[29][44] ;
wire \couts[29][43] ;
wire \couts[29][42] ;
wire \couts[29][41] ;
wire \couts[29][40] ;
wire \couts[29][39] ;
wire \couts[29][38] ;
wire \couts[29][37] ;
wire \couts[29][36] ;
wire \couts[29][35] ;
wire \couts[29][34] ;
wire \couts[29][33] ;
wire \couts[29][32] ;
wire \couts[29][31] ;
wire \couts[29][30] ;
wire \couts[29][29] ;
wire \couts[29][28] ;
wire \couts[29][27] ;
wire \couts[29][26] ;
wire \couts[29][25] ;
wire \couts[29][24] ;
wire \couts[29][23] ;
wire \couts[29][22] ;
wire \couts[29][21] ;
wire \couts[29][20] ;
wire \couts[29][19] ;
wire \couts[29][18] ;
wire \couts[29][17] ;
wire \couts[29][16] ;
wire \couts[29][15] ;
wire \couts[29][14] ;
wire \couts[29][13] ;
wire \couts[29][12] ;
wire \couts[29][11] ;
wire \couts[29][10] ;
wire \couts[29][9] ;
wire \sums[29][63] ;
wire \sums[29][62] ;
wire \sums[29][61] ;
wire \sums[29][60] ;
wire \sums[29][59] ;
wire \sums[29][58] ;
wire \sums[29][57] ;
wire \sums[29][56] ;
wire \sums[29][55] ;
wire \sums[29][54] ;
wire \sums[29][53] ;
wire \sums[29][52] ;
wire \sums[29][51] ;
wire \sums[29][50] ;
wire \sums[29][49] ;
wire \sums[29][48] ;
wire \sums[29][47] ;
wire \sums[29][46] ;
wire \sums[29][45] ;
wire \sums[29][44] ;
wire \sums[29][43] ;
wire \sums[29][42] ;
wire \sums[29][41] ;
wire \sums[29][40] ;
wire \sums[29][39] ;
wire \sums[29][38] ;
wire \sums[29][37] ;
wire \sums[29][36] ;
wire \sums[29][35] ;
wire \sums[29][34] ;
wire \sums[29][33] ;
wire \sums[29][32] ;
wire \sums[29][31] ;
wire \sums[29][30] ;
wire \sums[29][29] ;
wire \sums[29][28] ;
wire \sums[29][27] ;
wire \sums[29][26] ;
wire \sums[29][25] ;
wire \sums[29][24] ;
wire \sums[29][23] ;
wire \sums[29][22] ;
wire \sums[29][21] ;
wire \sums[29][20] ;
wire \sums[29][19] ;
wire \sums[29][18] ;
wire \sums[29][17] ;
wire \sums[29][16] ;
wire \sums[29][15] ;
wire \sums[29][14] ;
wire \sums[29][13] ;
wire \sums[29][12] ;
wire \sums[29][11] ;
wire \sums[29][10] ;
wire \sums[29][9] ;
wire \couts[30][63] ;
wire \couts[30][62] ;
wire \couts[30][61] ;
wire \couts[30][60] ;
wire \couts[30][59] ;
wire \couts[30][58] ;
wire \couts[30][57] ;
wire \couts[30][56] ;
wire \couts[30][55] ;
wire \couts[30][54] ;
wire \couts[30][53] ;
wire \couts[30][52] ;
wire \couts[30][51] ;
wire \couts[30][50] ;
wire \couts[30][49] ;
wire \couts[30][48] ;
wire \couts[30][47] ;
wire \couts[30][46] ;
wire \couts[30][45] ;
wire \couts[30][44] ;
wire \couts[30][43] ;
wire \couts[30][42] ;
wire \couts[30][41] ;
wire \couts[30][40] ;
wire \couts[30][39] ;
wire \couts[30][38] ;
wire \couts[30][37] ;
wire \couts[30][36] ;
wire \couts[30][35] ;
wire \couts[30][34] ;
wire \couts[30][33] ;
wire \couts[30][32] ;
wire \couts[30][31] ;
wire \couts[30][30] ;
wire \couts[30][29] ;
wire \couts[30][28] ;
wire \couts[30][27] ;
wire \couts[30][26] ;
wire \couts[30][25] ;
wire \couts[30][24] ;
wire \couts[30][23] ;
wire \couts[30][22] ;
wire \couts[30][21] ;
wire \couts[30][20] ;
wire \couts[30][19] ;
wire \couts[30][18] ;
wire \couts[30][17] ;
wire \couts[30][16] ;
wire \couts[30][15] ;
wire \couts[30][14] ;
wire \couts[30][13] ;
wire \couts[30][12] ;
wire \couts[30][11] ;
wire \couts[30][10] ;
wire \sums[30][63] ;
wire \sums[30][62] ;
wire \sums[30][61] ;
wire \sums[30][60] ;
wire \sums[30][59] ;
wire \sums[30][58] ;
wire \sums[30][57] ;
wire \sums[30][56] ;
wire \sums[30][55] ;
wire \sums[30][54] ;
wire \sums[30][53] ;
wire \sums[30][52] ;
wire \sums[30][51] ;
wire \sums[30][50] ;
wire \sums[30][49] ;
wire \sums[30][48] ;
wire \sums[30][47] ;
wire \sums[30][46] ;
wire \sums[30][45] ;
wire \sums[30][44] ;
wire \sums[30][43] ;
wire \sums[30][42] ;
wire \sums[30][41] ;
wire \sums[30][40] ;
wire \sums[30][39] ;
wire \sums[30][38] ;
wire \sums[30][37] ;
wire \sums[30][36] ;
wire \sums[30][35] ;
wire \sums[30][34] ;
wire \sums[30][33] ;
wire \sums[30][32] ;
wire \sums[30][31] ;
wire \sums[30][30] ;
wire \sums[30][29] ;
wire \sums[30][28] ;
wire \sums[30][27] ;
wire \sums[30][26] ;
wire \sums[30][25] ;
wire \sums[30][24] ;
wire \sums[30][23] ;
wire \sums[30][22] ;
wire \sums[30][21] ;
wire \sums[30][20] ;
wire \sums[30][19] ;
wire \sums[30][18] ;
wire \sums[30][17] ;
wire \sums[30][16] ;
wire \sums[30][15] ;
wire \sums[30][14] ;
wire \sums[30][13] ;
wire \sums[30][12] ;
wire \sums[30][11] ;
wire \sums[30][10] ;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire uc_57;
wire uc_58;
wire uc_59;
wire uc_60;
wire uc_61;
wire uc_62;
wire uc_63;
wire uc_64;
wire uc_65;
wire uc_66;
wire uc_67;
wire uc_68;
wire uc_69;
wire uc_70;
wire uc_71;
wire uc_72;
wire uc_73;
wire uc_74;
wire uc_75;
wire uc_76;
wire uc_77;
wire uc_78;
wire uc_79;
wire uc_80;
wire uc_81;
wire uc_82;
wire uc_83;
wire uc_84;
wire uc_85;
wire uc_86;
wire uc_87;
wire uc_88;
wire uc_89;
wire uc_90;
wire uc_91;
wire uc_92;
wire uc_93;
wire uc_94;
wire uc_95;
wire uc_96;
wire uc_97;
wire uc_98;
wire uc_99;
wire uc_100;
wire uc_101;
wire uc_102;
wire uc_103;
wire uc_104;
wire uc_105;
wire uc_106;
wire uc_107;
wire uc_108;
wire uc_109;
wire uc_110;
wire uc_111;
wire uc_112;
wire uc_113;
wire uc_114;
wire uc_115;
wire uc_116;
wire uc_117;
wire uc_118;
wire uc_119;
wire uc_120;
wire uc_121;
wire uc_122;
wire uc_123;
wire uc_124;
wire uc_125;
wire uc_126;
wire uc_127;
wire uc_128;
wire uc_129;
wire uc_130;
wire uc_131;
wire uc_132;
wire uc_133;
wire uc_134;
wire uc_135;
wire uc_136;
wire uc_137;
wire uc_138;
wire uc_139;
wire uc_140;
wire uc_141;
wire uc_142;
wire uc_143;
wire uc_144;
wire uc_145;
wire uc_146;
wire uc_147;
wire uc_148;
wire uc_149;
wire uc_150;
wire uc_151;
wire uc_152;
wire uc_153;
wire uc_154;
wire uc_155;
wire uc_156;
wire uc_157;
wire uc_158;
wire uc_159;
wire uc_160;
wire uc_161;
wire uc_162;
wire uc_163;
wire uc_164;
wire uc_165;
wire uc_166;
wire uc_167;
wire uc_168;
wire uc_169;
wire uc_170;
wire uc_171;
wire uc_172;
wire uc_173;
wire uc_174;
wire uc_175;
wire uc_176;
wire uc_177;
wire uc_178;
wire uc_179;
wire uc_180;
wire uc_181;
wire uc_182;
wire uc_183;
wire uc_184;
wire uc_185;
wire uc_186;
wire uc_187;
wire uc_188;
wire uc_189;
wire uc_190;
wire uc_191;
wire uc_192;
wire uc_193;
wire uc_194;
wire uc_195;
wire uc_196;
wire uc_197;
wire uc_198;
wire uc_199;
wire uc_200;
wire uc_201;
wire uc_202;
wire uc_203;
wire uc_204;
wire uc_205;
wire uc_206;
wire uc_207;
wire uc_208;
wire uc_209;
wire uc_210;
wire uc_211;
wire uc_212;
wire uc_213;
wire uc_214;
wire uc_215;
wire uc_216;
wire uc_217;
wire uc_218;
wire uc_219;
wire uc_220;
wire uc_221;
wire uc_222;
wire uc_223;
wire uc_224;
wire uc_225;
wire uc_226;
wire uc_227;
wire uc_228;
wire uc_229;
wire uc_230;
wire uc_231;
wire uc_232;
wire uc_233;
wire uc_234;
wire uc_235;
wire uc_236;
wire uc_237;
wire uc_238;
wire uc_239;
wire uc_240;
wire uc_241;
wire uc_242;
wire uc_243;
wire uc_244;
wire uc_245;
wire uc_246;
wire uc_247;
wire uc_248;
wire uc_249;
wire uc_250;
wire uc_251;
wire uc_252;
wire uc_253;
wire uc_254;
wire uc_255;
wire uc_256;
wire uc_257;
wire uc_258;
wire uc_259;
wire uc_260;
wire uc_261;
wire uc_262;
wire uc_263;
wire uc_264;
wire uc_265;
wire uc_266;
wire uc_267;
wire uc_268;
wire uc_269;
wire uc_270;
wire uc_271;
wire uc_272;
wire uc_273;
wire uc_274;
wire uc_275;
wire uc_276;
wire uc_277;
wire uc_278;
wire uc_279;
wire uc_280;
wire uc_281;
wire uc_282;
wire uc_283;
wire uc_284;
wire uc_285;
wire uc_286;
wire uc_287;
wire uc_288;
wire uc_289;
wire uc_290;
wire uc_291;
wire uc_292;
wire uc_293;
wire uc_294;
wire uc_295;
wire uc_296;
wire uc_297;
wire uc_298;
wire uc_299;
wire uc_300;
wire uc_301;
wire uc_302;
wire uc_303;
wire uc_304;
wire uc_305;
wire uc_306;
wire uc_307;
wire uc_308;
wire uc_309;
wire uc_310;
wire uc_311;
wire uc_312;
wire uc_313;
wire uc_314;
wire uc_315;
wire uc_316;
wire uc_317;
wire uc_318;
wire uc_319;
wire uc_320;
wire uc_321;
wire uc_322;
wire uc_323;
wire uc_324;
wire uc_325;
wire uc_326;
wire uc_327;
wire uc_328;
wire uc_329;
wire uc_330;
wire uc_331;
wire uc_332;
wire uc_333;
wire uc_334;
wire uc_335;
wire uc_336;
wire uc_337;
wire uc_338;
wire uc_339;
wire uc_340;
wire uc_341;
wire uc_342;
wire uc_343;
wire uc_344;
wire uc_345;
wire uc_346;
wire uc_347;
wire uc_348;
wire uc_349;
wire uc_350;
wire uc_351;
wire uc_352;
wire uc_353;
wire uc_354;
wire uc_355;
wire uc_356;
wire uc_357;
wire uc_358;
wire uc_359;
wire uc_360;
wire uc_361;
wire uc_362;
wire uc_363;
wire uc_364;
wire uc_365;
wire uc_366;
wire uc_367;
wire uc_368;
wire uc_369;
wire uc_370;
wire uc_371;
wire uc_372;
wire uc_373;
wire uc_374;
wire uc_375;
wire uc_376;
wire uc_377;
wire uc_378;
wire uc_379;
wire uc_380;
wire uc_381;
wire uc_382;
wire uc_383;
wire uc_384;
wire uc_385;
wire uc_386;
wire uc_387;
wire uc_388;
wire uc_389;
wire uc_390;
wire uc_391;
wire uc_392;
wire uc_393;
wire uc_394;
wire uc_395;
wire uc_396;
wire uc_397;
wire uc_398;
wire uc_399;
wire uc_400;
wire uc_401;
wire uc_402;
wire uc_403;
wire uc_404;
wire uc_405;
wire uc_406;
wire uc_407;
wire uc_408;
wire uc_409;
wire uc_410;
wire uc_411;
wire uc_412;
wire uc_413;
wire uc_414;
wire uc_415;
wire uc_416;
wire uc_417;
wire uc_418;
wire uc_419;
wire uc_420;
wire uc_421;
wire uc_422;
wire uc_423;
wire uc_424;
wire uc_425;
wire uc_426;
wire uc_427;
wire uc_428;
wire uc_429;
wire uc_430;
wire uc_431;
wire uc_432;
wire uc_433;
wire uc_434;
wire uc_435;
wire uc_436;
wire uc_437;
wire uc_438;
wire uc_439;
wire uc_440;
wire uc_441;
wire uc_442;
wire uc_443;
wire uc_444;
wire uc_445;
wire uc_446;
wire uc_447;
wire uc_448;
wire uc_449;
wire uc_450;
wire uc_451;
wire uc_452;
wire uc_453;
wire uc_454;
wire uc_455;
wire uc_456;
wire uc_457;
wire uc_458;
wire uc_459;
wire uc_460;
wire uc_461;
wire uc_462;
wire uc_463;
wire uc_464;
wire uc_465;
wire uc_466;
wire uc_467;
wire uc_468;
wire uc_469;
wire uc_470;
wire uc_471;
wire uc_472;
wire uc_473;
wire uc_474;
wire uc_475;
wire uc_476;
wire uc_477;
wire uc_478;
wire uc_479;
wire uc_480;
wire uc_481;
wire uc_482;
wire uc_483;
wire uc_484;
wire uc_485;
wire uc_486;
wire uc_487;
wire uc_488;
wire uc_489;
wire uc_490;
wire uc_491;
wire uc_492;
wire uc_493;
wire uc_494;
wire uc_495;
wire uc_496;
wire uc_497;
wire uc_498;
wire uc_499;
wire uc_500;
wire uc_501;
wire uc_502;
wire uc_503;
wire uc_504;
wire uc_505;
wire uc_506;
wire uc_507;
wire uc_508;
wire uc_509;
wire uc_510;
wire uc_511;
wire uc_512;
wire uc_513;
wire uc_514;
wire uc_515;
wire uc_516;
wire uc_517;
wire uc_518;
wire uc_519;
wire uc_520;
wire uc_521;
wire uc_522;
wire uc_523;
wire uc_524;
wire uc_525;
wire uc_526;
wire uc_527;
wire uc_528;
wire uc_529;
wire uc_530;
wire uc_531;
wire uc_532;
wire uc_533;
wire uc_534;
wire uc_535;
wire uc_536;
wire uc_537;
wire uc_538;
wire uc_539;
wire uc_540;
wire uc_541;
wire uc_542;
wire uc_543;
wire uc_544;
wire uc_545;
wire uc_546;
wire uc_547;
wire uc_548;
wire uc_549;
wire uc_550;
wire uc_551;
wire uc_552;
wire uc_553;
wire uc_554;
wire uc_555;
wire uc_556;
wire uc_557;
wire uc_558;
wire uc_559;
wire uc_560;
wire uc_561;
wire uc_562;
wire uc_563;
wire uc_564;
wire uc_565;
wire uc_566;
wire uc_567;
wire uc_568;
wire uc_569;
wire uc_570;
wire uc_571;
wire uc_572;
wire uc_573;
wire uc_574;
wire uc_575;
wire uc_576;
wire uc_577;
wire uc_578;
wire uc_579;
wire uc_580;
wire uc_581;
wire uc_582;
wire uc_583;
wire uc_584;
wire uc_585;
wire uc_586;
wire uc_587;
wire uc_588;
wire uc_589;
wire uc_590;
wire uc_591;
wire uc_592;
wire uc_593;
wire uc_594;
wire uc_595;
wire uc_596;
wire uc_597;
wire uc_598;
wire uc_599;
wire uc_600;
wire uc_601;
wire uc_602;
wire uc_603;
wire uc_604;
wire uc_605;
wire uc_606;
wire uc_607;
wire uc_608;
wire uc_609;
wire uc_610;
wire uc_611;
wire uc_612;
wire uc_613;
wire uc_614;
wire uc_615;
wire uc_616;
wire uc_617;
wire uc_618;
wire uc_619;
wire uc_620;
wire uc_621;
wire uc_622;
wire uc_623;
wire uc_624;
wire uc_625;
wire uc_626;
wire uc_627;
wire uc_628;
wire uc_629;
wire uc_630;
wire uc_631;
wire uc_632;
wire uc_633;
wire uc_634;
wire uc_635;
wire uc_636;
wire uc_637;
wire uc_638;
wire uc_639;
wire uc_640;
wire uc_641;
wire uc_642;
wire uc_643;
wire uc_644;
wire uc_645;
wire uc_646;
wire uc_647;
wire uc_648;
wire uc_649;
wire uc_650;
wire uc_651;
wire uc_652;
wire uc_653;
wire uc_654;
wire uc_655;
wire uc_656;
wire uc_657;
wire uc_658;
wire uc_659;
wire uc_660;
wire uc_661;
wire uc_662;
wire uc_663;
wire uc_664;
wire uc_665;
wire uc_666;
wire uc_667;
wire uc_668;
wire uc_669;
wire uc_670;
wire uc_671;
wire uc_672;
wire uc_673;
wire uc_674;
wire uc_675;
wire uc_676;
wire uc_677;
wire uc_678;
wire uc_679;
wire uc_680;
wire uc_681;
wire uc_682;
wire uc_683;
wire uc_684;
wire uc_685;
wire uc_686;
wire uc_687;
wire uc_688;
wire uc_689;
wire uc_690;
wire uc_691;
wire uc_692;
wire uc_693;
wire uc_694;
wire uc_695;
wire uc_696;
wire uc_697;
wire uc_698;
wire uc_699;
wire uc_700;
wire uc_701;
wire uc_702;
wire uc_703;
wire uc_704;
wire uc_705;
wire uc_706;
wire uc_707;
wire uc_708;
wire uc_709;
wire uc_710;
wire uc_711;
wire uc_712;
wire uc_713;
wire uc_714;
wire uc_715;
wire uc_716;
wire uc_717;
wire uc_718;
wire uc_719;
wire uc_720;
wire uc_721;
wire uc_722;
wire uc_723;
wire uc_724;
wire uc_725;
wire uc_726;
wire uc_727;
wire uc_728;
wire uc_729;
wire uc_730;
wire uc_731;
wire uc_732;
wire uc_733;
wire uc_734;
wire uc_735;
wire uc_736;
wire uc_737;
wire uc_738;
wire uc_739;
wire uc_740;
wire uc_741;
wire uc_742;
wire uc_743;
wire uc_744;
wire uc_745;
wire uc_746;
wire uc_747;
wire uc_748;
wire uc_749;
wire uc_750;
wire uc_751;
wire uc_752;
wire uc_753;
wire uc_754;
wire uc_755;
wire uc_756;
wire uc_757;
wire uc_758;
wire uc_759;
wire uc_760;
wire uc_761;
wire uc_762;
wire uc_763;
wire uc_764;
wire uc_765;
wire uc_766;
wire uc_767;
wire uc_768;
wire uc_769;
wire uc_770;
wire uc_771;
wire uc_772;
wire uc_773;
wire uc_774;
wire uc_775;
wire uc_776;
wire uc_777;
wire uc_778;
wire uc_779;
wire uc_780;
wire uc_781;
wire uc_782;
wire uc_783;
wire uc_784;
wire uc_785;
wire uc_786;
wire uc_787;
wire uc_788;
wire uc_789;
wire uc_790;
wire uc_791;
wire uc_792;
wire uc_793;
wire uc_794;
wire uc_795;
wire uc_796;
wire uc_797;
wire uc_798;
wire uc_799;
wire uc_800;
wire uc_801;
wire uc_802;
wire uc_803;
wire uc_804;
wire uc_805;
wire uc_806;
wire uc_807;
wire uc_808;
wire uc_809;
wire uc_810;
wire uc_811;
wire uc_812;
wire uc_813;
wire uc_814;
wire uc_815;
wire uc_816;
wire uc_817;
wire uc_818;
wire uc_819;
wire uc_820;
wire uc_821;
wire uc_822;
wire uc_823;
wire uc_824;
wire uc_825;
wire uc_826;
wire uc_827;
wire uc_828;
wire uc_829;
wire uc_830;
wire uc_831;
wire uc_832;
wire uc_833;
wire uc_834;
wire uc_835;
wire uc_836;
wire uc_837;
wire uc_838;
wire uc_839;
wire uc_840;
wire uc_841;
wire uc_842;
wire uc_843;
wire uc_844;
wire uc_845;
wire uc_846;
wire uc_847;
wire uc_848;
wire uc_849;
wire uc_850;
wire uc_851;
wire uc_852;
wire uc_853;
wire uc_854;
wire uc_855;
wire uc_856;
wire uc_857;
wire uc_858;
wire uc_859;
wire uc_860;
wire uc_861;
wire uc_862;
wire uc_863;
wire uc_864;
wire uc_865;
wire uc_866;
wire uc_867;
wire uc_868;
wire uc_869;
wire uc_870;
wire uc_871;
wire uc_872;
wire uc_873;
wire uc_874;
wire uc_875;
wire uc_876;
wire uc_877;
wire uc_878;
wire uc_879;
wire uc_880;
wire uc_881;
wire uc_882;
wire uc_883;
wire uc_884;
wire uc_885;
wire uc_886;
wire uc_887;
wire uc_888;
wire uc_889;
wire uc_890;
wire uc_891;
wire uc_892;
wire uc_893;
wire uc_894;
wire uc_895;
wire uc_896;
wire uc_897;
wire uc_898;
wire uc_899;
wire uc_900;
wire uc_901;
wire uc_902;
wire uc_903;
wire uc_904;
wire uc_905;
wire uc_906;
wire uc_907;
wire uc_908;
wire uc_909;
wire uc_910;
wire uc_911;
wire uc_912;
wire uc_913;
wire uc_914;
wire uc_915;
wire uc_916;
wire uc_917;
wire uc_918;
wire uc_919;
wire uc_920;
wire uc_921;
wire uc_922;
wire uc_923;
wire uc_924;
wire uc_925;
wire uc_926;
wire uc_927;
wire uc_928;
wire uc_929;
wire uc_930;
wire uc_931;
wire uc_932;
wire uc_933;
wire uc_934;
wire uc_935;
wire uc_936;
wire uc_937;
wire uc_938;
wire uc_939;
wire uc_940;
wire uc_941;
wire uc_942;
wire uc_943;
wire uc_944;
wire uc_945;
wire uc_946;
wire uc_947;
wire uc_948;
wire uc_949;
wire uc_950;
wire uc_951;
wire uc_952;
wire uc_953;
wire uc_954;
wire uc_955;
wire uc_956;
wire uc_957;
wire uc_958;
wire uc_959;
wire uc_960;
wire uc_961;
wire uc_962;
wire uc_963;
wire uc_964;
wire uc_965;
wire uc_966;
wire uc_967;
wire uc_968;
wire uc_969;
wire uc_970;
wire uc_971;
wire uc_972;
wire uc_973;
wire uc_974;
wire uc_975;
wire uc_976;
wire uc_977;
wire uc_978;
wire uc_979;
wire uc_980;
wire uc_981;
wire uc_982;
wire uc_983;
wire uc_984;
wire uc_985;
wire uc_986;
wire uc_987;
wire uc_988;
wire uc_989;
wire uc_990;
wire uc_991;
wire uc_992;
wire uc_993;
wire uc_994;
wire uc_995;
wire uc_996;
wire uc_997;
wire uc_998;
wire uc_999;
wire uc_1000;
wire uc_1001;
wire uc_1002;
wire uc_1003;
wire uc_1004;
wire uc_1005;
wire uc_1006;
wire uc_1007;
wire uc_1008;
wire uc_1009;
wire uc_1010;
wire uc_1011;
wire uc_1012;
wire uc_1013;
wire uc_1014;
wire uc_1015;
wire uc_1016;
wire uc_1017;
wire uc_1018;
wire uc_1019;
wire uc_1020;
wire uc_1021;
wire uc_1022;
wire uc_1023;
wire uc_1024;
wire uc_1025;
wire uc_1026;
wire uc_1027;
wire uc_1028;
wire uc_1029;
wire uc_1030;
wire uc_1031;
wire uc_1032;
wire uc_1033;
wire uc_1034;
wire uc_1035;
wire uc_1036;
wire uc_1037;
wire uc_1038;
wire uc_1039;
wire uc_1040;
wire uc_1041;
wire uc_1042;
wire uc_1043;
wire uc_1044;
wire uc_1045;
wire uc_1046;
wire uc_1047;
wire uc_1048;
wire uc_1049;
wire uc_1050;
wire uc_1051;
wire uc_1052;
wire uc_1053;
wire uc_1054;
wire uc_1055;
wire uc_1056;
wire uc_1057;
wire uc_1058;
wire uc_1059;
wire uc_1060;
wire uc_1061;
wire uc_1062;
wire uc_1063;
wire uc_1064;
wire uc_1065;
wire uc_1066;
wire uc_1067;
wire uc_1068;
wire uc_1069;
wire uc_1070;
wire uc_1071;
wire uc_1072;
wire uc_1073;
wire uc_1074;
wire uc_1075;
wire uc_1076;
wire uc_1077;
wire uc_1078;
wire uc_1079;
wire uc_1080;
wire uc_1081;
wire uc_1082;
wire uc_1083;
wire uc_1084;
wire uc_1085;
wire uc_1086;
wire uc_1087;
wire uc_1088;
wire uc_1089;
wire uc_1090;
wire uc_1091;
wire uc_1092;
wire uc_1093;
wire uc_1094;
wire uc_1095;
wire uc_1096;
wire uc_1097;
wire uc_1098;
wire uc_1099;
wire uc_1100;
wire uc_1101;
wire uc_1102;
wire uc_1103;
wire uc_1104;
wire uc_1105;
wire uc_1106;
wire uc_1107;
wire uc_1108;
wire uc_1109;
wire uc_1110;
wire uc_1111;
wire uc_1112;
wire uc_1113;
wire uc_1114;
wire uc_1115;
wire uc_1116;
wire uc_1117;
wire uc_1118;
wire uc_1119;
wire uc_1120;
wire uc_1121;
wire uc_1122;
wire uc_1123;
wire uc_1124;
wire uc_1125;
wire uc_1126;
wire uc_1127;
wire uc_1128;
wire uc_1129;
wire uc_1130;
wire uc_1131;
wire uc_1132;
wire uc_1133;
wire uc_1134;
wire uc_1135;
wire uc_1136;
wire uc_1137;
wire uc_1138;
wire uc_1139;
wire uc_1140;
wire uc_1141;
wire uc_1142;
wire uc_1143;
wire uc_1144;
wire uc_1145;
wire uc_1146;
wire uc_1147;
wire uc_1148;
wire uc_1149;
wire uc_1150;
wire uc_1151;
wire uc_1152;
wire uc_1153;
wire uc_1154;
wire uc_1155;
wire uc_1156;
wire uc_1157;
wire uc_1158;
wire uc_1159;
wire uc_1160;
wire uc_1161;
wire uc_1162;
wire uc_1163;
wire uc_1164;
wire uc_1165;
wire uc_1166;
wire uc_1167;
wire uc_1168;
wire uc_1169;
wire uc_1170;
wire uc_1171;
wire uc_1172;
wire uc_1173;
wire uc_1174;
wire uc_1175;
wire uc_1176;
wire uc_1177;
wire uc_1178;
wire uc_1179;
wire uc_1180;
wire uc_1181;
wire uc_1182;
wire uc_1183;
wire uc_1184;
wire uc_1185;
wire uc_1186;
wire uc_1187;
wire uc_1188;
wire uc_1189;
wire uc_1190;
wire uc_1191;
wire uc_1192;
wire uc_1193;
wire uc_1194;
wire uc_1195;
wire uc_1196;
wire uc_1197;
wire uc_1198;
wire uc_1199;
wire uc_1200;
wire uc_1201;
wire uc_1202;
wire uc_1203;
wire uc_1204;
wire uc_1205;
wire uc_1206;
wire uc_1207;
wire uc_1208;
wire uc_1209;
wire uc_1210;
wire uc_1211;
wire uc_1212;
wire uc_1213;
wire uc_1214;
wire uc_1215;
wire uc_1216;
wire uc_1217;
wire uc_1218;
wire uc_1219;
wire uc_1220;
wire uc_1221;
wire uc_1222;
wire uc_1223;
wire uc_1224;
wire uc_1225;
wire uc_1226;
wire uc_1227;
wire uc_1228;
wire uc_1229;
wire uc_1230;
wire uc_1231;
wire uc_1232;
wire uc_1233;
wire uc_1234;
wire uc_1235;
wire uc_1236;
wire uc_1237;
wire uc_1238;
wire uc_1239;
wire uc_1240;
wire uc_1241;
wire uc_1242;
wire uc_1243;
wire uc_1244;
wire uc_1245;
wire uc_1246;
wire uc_1247;
wire uc_1248;
wire uc_1249;
wire uc_1250;
wire uc_1251;
wire uc_1252;
wire uc_1253;
wire uc_1254;
wire uc_1255;
wire uc_1256;
wire uc_1257;
wire uc_1258;
wire uc_1259;
wire uc_1260;
wire uc_1261;
wire uc_1262;
wire uc_1263;
wire uc_1264;
wire uc_1265;
wire uc_1266;
wire uc_1267;
wire uc_1268;
wire uc_1269;
wire uc_1270;
wire uc_1271;
wire uc_1272;
wire uc_1273;
wire uc_1274;
wire uc_1275;
wire uc_1276;
wire uc_1277;
wire uc_1278;
wire uc_1279;
wire uc_1280;
wire uc_1281;
wire uc_1282;
wire uc_1283;
wire uc_1284;
wire uc_1285;
wire uc_1286;
wire uc_1287;
wire uc_1288;
wire uc_1289;
wire uc_1290;
wire uc_1291;
wire uc_1292;
wire uc_1293;
wire uc_1294;
wire uc_1295;
wire uc_1296;
wire uc_1297;
wire uc_1298;
wire uc_1299;
wire uc_1300;
wire uc_1301;
wire uc_1302;
wire uc_1303;
wire uc_1304;
wire uc_1305;
wire uc_1306;
wire uc_1307;
wire uc_1308;
wire uc_1309;
wire uc_1310;
wire uc_1311;
wire uc_1312;
wire uc_1313;
wire uc_1314;
wire uc_1315;
wire uc_1316;
wire uc_1317;
wire uc_1318;
wire uc_1319;
wire uc_1320;
wire uc_1321;
wire uc_1322;
wire uc_1323;
wire uc_1324;
wire uc_1325;
wire uc_1326;
wire uc_1327;
wire uc_1328;
wire uc_1329;
wire uc_1330;
wire uc_1331;
wire uc_1332;
wire uc_1333;
wire uc_1334;
wire uc_1335;
wire uc_1336;
wire uc_1337;
wire uc_1338;
wire uc_1339;
wire uc_1340;
wire uc_1341;
wire uc_1342;
wire uc_1343;
wire uc_1344;
wire uc_1345;
wire uc_1346;
wire uc_1347;
wire uc_1348;
wire uc_1349;
wire uc_1350;
wire uc_1351;
wire uc_1352;
wire uc_1353;
wire uc_1354;
wire uc_1355;
wire uc_1356;
wire uc_1357;
wire uc_1358;
wire uc_1359;
wire uc_1360;
wire uc_1361;
wire uc_1362;
wire uc_1363;
wire uc_1364;
wire uc_1365;
wire uc_1366;
wire uc_1367;
wire uc_1368;
wire uc_1369;
wire uc_1370;
wire uc_1371;
wire uc_1372;
wire uc_1373;
wire uc_1374;
wire uc_1375;
wire uc_1376;
wire uc_1377;
wire uc_1378;
wire uc_1379;
wire uc_1380;
wire uc_1381;
wire uc_1382;
wire uc_1383;
wire uc_1384;
wire uc_1385;
wire uc_1386;
wire uc_1387;
wire uc_1388;
wire uc_1389;
wire uc_1390;
wire uc_1391;
wire uc_1392;
wire uc_1393;
wire uc_1394;
wire uc_1395;
wire uc_1396;
wire uc_1397;
wire uc_1398;
wire uc_1399;
wire uc_1400;
wire uc_1401;
wire uc_1402;
wire uc_1403;
wire uc_1404;
wire uc_1405;
wire uc_1406;
wire uc_1407;
wire uc_1408;
wire uc_1409;
wire uc_1410;
wire uc_1411;
wire uc_1412;
wire uc_1413;
wire uc_1414;
wire uc_1415;
wire uc_1416;
wire uc_1417;
wire uc_1418;
wire uc_1419;
wire uc_1420;
wire uc_1421;
wire uc_1422;
wire uc_1423;
wire uc_1424;
wire uc_1425;
wire uc_1426;
wire uc_1427;
wire uc_1428;
wire uc_1429;
wire uc_1430;
wire uc_1431;
wire uc_1432;
wire uc_1433;
wire uc_1434;
wire uc_1435;
wire uc_1436;
wire uc_1437;
wire uc_1438;
wire uc_1439;
wire uc_1440;
wire uc_1441;
wire uc_1442;
wire uc_1443;
wire uc_1444;
wire uc_1445;
wire uc_1446;
wire uc_1447;
wire uc_1448;
wire uc_1449;
wire uc_1450;
wire uc_1451;
wire uc_1452;
wire uc_1453;
wire uc_1454;
wire uc_1455;
wire uc_1456;
wire uc_1457;
wire uc_1458;
wire uc_1459;
wire uc_1460;
wire uc_1461;
wire uc_1462;
wire uc_1463;
wire uc_1464;
wire uc_1465;
wire uc_1466;
wire uc_1467;
wire uc_1468;
wire uc_1469;
wire uc_1470;
wire uc_1471;
wire uc_1472;
wire uc_1473;
wire uc_1474;
wire uc_1475;
wire uc_1476;
wire uc_1477;
wire uc_1478;
wire uc_1479;
wire uc_1480;
wire uc_1481;
wire uc_1482;
wire uc_1483;
wire uc_1484;
wire uc_1485;
wire uc_1486;
wire uc_1487;
wire uc_1488;
wire uc_1489;
wire uc_1490;
wire uc_1491;
wire uc_1492;
wire uc_1493;
wire uc_1494;
wire uc_1495;
wire uc_1496;
wire uc_1497;
wire uc_1498;
wire uc_1499;
wire uc_1500;
wire uc_1501;
wire uc_1502;
wire uc_1503;
wire uc_1504;
wire uc_1505;
wire uc_1506;
wire uc_1507;
wire uc_1508;
wire uc_1509;
wire uc_1510;
wire uc_1511;
wire uc_1512;
wire uc_1513;
wire uc_1514;
wire uc_1515;
wire uc_1516;
wire uc_1517;
wire uc_1518;
wire uc_1519;
wire uc_1520;
wire uc_1521;
wire uc_1522;
wire uc_1523;
wire uc_1524;
wire uc_1525;
wire uc_1526;
wire uc_1527;
wire uc_1528;
wire uc_1529;
wire uc_1530;
wire uc_1531;
wire uc_1532;
wire uc_1533;
wire uc_1534;
wire uc_1535;
wire uc_1536;
wire uc_1537;
wire uc_1538;
wire uc_1539;
wire uc_1540;
wire uc_1541;
wire uc_1542;
wire uc_1543;
wire uc_1544;
wire uc_1545;
wire uc_1546;
wire uc_1547;
wire uc_1548;
wire uc_1549;
wire uc_1550;
wire uc_1551;
wire uc_1552;
wire uc_1553;
wire uc_1554;
wire uc_1555;
wire uc_1556;
wire uc_1557;
wire uc_1558;
wire uc_1559;
wire uc_1560;
wire uc_1561;
wire uc_1562;
wire uc_1563;
wire uc_1564;
wire uc_1565;
wire uc_1566;
wire uc_1567;
wire uc_1568;
wire uc_1569;
wire uc_1570;
wire uc_1571;
wire uc_1572;
wire uc_1573;
wire uc_1574;
wire uc_1575;
wire uc_1576;
wire uc_1577;
wire uc_1578;
wire uc_1579;
wire uc_1580;
wire uc_1581;
wire uc_1582;
wire uc_1583;
wire uc_1584;
wire uc_1585;
wire uc_1586;
wire uc_1587;
wire uc_1588;
wire uc_1589;
wire uc_1590;
wire uc_1591;
wire uc_1592;
wire uc_1593;
wire uc_1594;
wire uc_1595;
wire uc_1596;
wire uc_1597;
wire uc_1598;
wire uc_1599;
wire uc_1600;
wire uc_1601;
wire uc_1602;
wire uc_1603;
wire uc_1604;
wire uc_1605;
wire uc_1606;
wire uc_1607;
wire uc_1608;
wire uc_1609;
wire uc_1610;
wire uc_1611;
wire uc_1612;
wire uc_1613;
wire uc_1614;
wire uc_1615;
wire uc_1616;
wire uc_1617;
wire uc_1618;
wire uc_1619;
wire uc_1620;
wire uc_1621;
wire uc_1622;
wire uc_1623;
wire uc_1624;
wire uc_1625;
wire uc_1626;
wire uc_1627;
wire uc_1628;
wire uc_1629;
wire uc_1630;
wire uc_1631;
wire uc_1632;
wire uc_1633;
wire uc_1634;
wire uc_1635;
wire uc_1636;
wire uc_1637;
wire uc_1638;
wire uc_1639;
wire uc_1640;
wire uc_1641;
wire uc_1642;
wire uc_1643;
wire uc_1644;
wire uc_1645;
wire uc_1646;
wire uc_1647;
wire uc_1648;
wire uc_1649;
wire uc_1650;
wire uc_1651;
wire uc_1652;
wire uc_1653;
wire uc_1654;
wire uc_1655;
wire uc_1656;
wire uc_1657;
wire uc_1658;
wire uc_1659;
wire uc_1660;
wire uc_1661;
wire uc_1662;
wire uc_1663;
wire uc_1664;
wire uc_1665;
wire uc_1666;
wire uc_1667;
wire uc_1668;
wire uc_1669;
wire uc_1670;
wire uc_1671;
wire uc_1672;
wire uc_1673;
wire uc_1674;
wire uc_1675;
wire uc_1676;
wire uc_1677;
wire uc_1678;
wire uc_1679;
wire uc_1680;
wire uc_1681;
wire uc_1682;
wire uc_1683;
wire uc_1684;
wire uc_1685;
wire uc_1686;
wire uc_1687;
wire uc_1688;
wire uc_1689;
wire uc_1690;
wire uc_1691;
wire uc_1692;
wire uc_1693;
wire uc_1694;
wire uc_1695;
wire uc_1696;
wire uc_1697;
wire uc_1698;
wire uc_1699;
wire uc_1700;
wire uc_1701;
wire uc_1702;
wire uc_1703;
wire uc_1704;
wire uc_1705;
wire uc_1706;
wire uc_1707;
wire uc_1708;
wire uc_1709;
wire uc_1710;
wire uc_1711;
wire uc_1712;
wire uc_1713;
wire uc_1714;
wire uc_1715;
wire uc_1716;
wire uc_1717;
wire uc_1718;
wire uc_1719;
wire uc_1720;
wire uc_1721;
wire uc_1722;
wire uc_1723;
wire uc_1724;
wire uc_1725;
wire uc_1726;
wire uc_1727;
wire uc_1728;
wire uc_1729;
wire uc_1730;
wire uc_1731;
wire uc_1732;
wire uc_1733;
wire uc_1734;
wire uc_1735;
wire uc_1736;
wire uc_1737;
wire uc_1738;
wire uc_1739;
wire uc_1740;
wire uc_1741;
wire uc_1742;
wire uc_1743;
wire uc_1744;
wire uc_1745;
wire uc_1746;
wire uc_1747;
wire uc_1748;
wire uc_1749;
wire uc_1750;
wire uc_1751;
wire uc_1752;
wire uc_1753;
wire uc_1754;
wire uc_1755;
wire uc_1756;
wire uc_1757;
wire uc_1758;
wire uc_1759;
wire uc_1760;
wire uc_1761;
wire uc_1762;
wire uc_1763;
wire uc_1764;
wire uc_1765;
wire uc_1766;
wire uc_1767;
wire uc_1768;
wire uc_1769;
wire uc_1770;
wire uc_1771;
wire uc_1772;
wire uc_1773;
wire uc_1774;
wire uc_1775;
wire uc_1776;
wire uc_1777;
wire uc_1778;
wire uc_1779;
wire uc_1780;
wire uc_1781;
wire uc_1782;
wire uc_1783;
wire uc_1784;
wire uc_1785;
wire uc_1786;
wire uc_1787;
wire uc_1788;
wire uc_1789;
wire uc_1790;
wire uc_1791;
wire uc_1792;
wire uc_1793;
wire uc_1794;
wire uc_1795;
wire uc_1796;
wire uc_1797;
wire uc_1798;
wire uc_1799;
wire uc_1800;
wire uc_1801;
wire uc_1802;
wire uc_1803;
wire uc_1804;
wire uc_1805;
wire uc_1806;
wire uc_1807;
wire uc_1808;
wire uc_1809;
wire uc_1810;
wire uc_1811;
wire uc_1812;
wire uc_1813;
wire uc_1814;
wire uc_1815;
wire uc_1816;
wire uc_1817;
wire uc_1818;
wire uc_1819;
wire uc_1820;
wire uc_1821;
wire uc_1822;
wire uc_1823;
wire uc_1824;
wire uc_1825;
wire uc_1826;
wire uc_1827;
wire uc_1828;
wire uc_1829;
wire uc_1830;
wire uc_1831;
wire uc_1832;
wire uc_1833;
wire uc_1834;
wire uc_1835;
wire uc_1836;
wire uc_1837;
wire uc_1838;
wire uc_1839;
wire uc_1840;
wire uc_1841;
wire uc_1842;
wire uc_1843;
wire uc_1844;
wire uc_1845;
wire uc_1846;
wire uc_1847;
wire uc_1848;
wire uc_1849;
wire uc_1850;
wire uc_1851;
wire uc_1852;
wire uc_1853;
wire uc_1854;
wire uc_1855;
wire uc_1856;
wire uc_1857;
wire uc_1858;
wire uc_1859;
wire uc_1860;
wire uc_1861;
wire uc_1862;
wire uc_1863;
wire uc_1864;
wire uc_1865;
wire uc_1866;
wire uc_1867;
wire uc_1868;
wire uc_1869;
wire uc_1870;
wire uc_1871;
wire uc_1872;
wire uc_1873;
wire uc_1874;
wire uc_1875;
wire uc_1876;
wire uc_1877;
wire uc_1878;
wire uc_1879;
wire uc_1880;
wire uc_1881;
wire uc_1882;
wire uc_1883;
wire uc_1884;
wire uc_1885;
wire uc_1886;
wire uc_1887;
wire uc_1888;
wire uc_1889;
wire uc_1890;
wire uc_1891;
wire uc_1892;
wire uc_1893;
wire uc_1894;
wire uc_1895;
wire uc_1896;
wire uc_1897;
wire uc_1898;
wire uc_1899;
wire uc_1900;
wire uc_1901;
wire uc_1902;
wire uc_1903;
wire uc_1904;
wire uc_1905;
wire uc_1906;
wire uc_1907;
wire uc_1908;
wire uc_1909;
wire uc_1910;
wire uc_1911;
wire uc_1912;
wire uc_1913;
wire uc_1914;
wire uc_1915;
wire uc_1916;
wire uc_1917;
wire uc_1918;
wire uc_1919;
wire uc_1920;
wire uc_1921;
wire uc_1922;
wire uc_1923;
wire uc_1924;
wire uc_1925;
wire uc_1926;
wire uc_1927;
wire uc_1928;
wire uc_1929;
wire uc_1930;
wire uc_1931;
wire uc_1932;
wire uc_1933;
wire uc_1934;
wire uc_1935;
wire uc_1936;
wire uc_1937;
wire uc_1938;
wire uc_1939;
wire uc_1940;
wire uc_1941;
wire uc_1942;
wire uc_1943;
wire uc_1944;
wire uc_1945;
wire uc_1946;
wire uc_1947;
wire uc_1948;
wire uc_1949;
wire uc_1950;
wire uc_1951;
wire uc_1952;
wire uc_1953;
wire uc_1954;
wire uc_1955;
wire uc_1956;
wire uc_1957;
wire uc_1958;
wire uc_1959;
wire uc_1960;
wire uc_1961;
wire uc_1962;
wire uc_1963;
wire uc_1964;
wire uc_1965;
wire uc_1966;
wire uc_1967;
wire uc_1968;
wire uc_1969;
wire uc_1970;
wire uc_1971;
wire uc_1972;
wire uc_1973;
wire uc_1974;
wire uc_1975;
wire uc_1976;
wire uc_1977;
wire uc_1978;
wire uc_1979;
wire uc_1980;
wire uc_1981;
wire uc_1982;
wire uc_1983;
wire uc_1984;
wire uc_1985;
wire uc_1986;
wire uc_1987;
wire uc_1988;
wire uc_1989;
wire uc_1990;
wire uc_1991;
wire uc_1992;
wire uc_1993;
wire uc_1994;
wire uc_1995;
wire uc_1996;
wire uc_1997;
wire uc_1998;
wire uc_1999;
wire uc_2000;
wire uc_2001;
wire uc_2002;
wire uc_2003;
wire uc_2004;
wire uc_2005;
wire uc_2006;
wire uc_2007;
wire uc_2008;
wire uc_2009;
wire uc_2010;
wire uc_2011;
wire uc_2012;
wire uc_2013;
wire uc_2014;
wire uc_2015;
wire uc_2016;
wire uc_2017;
wire uc_2018;
wire uc_2019;
wire uc_2020;
wire uc_2021;
wire uc_2022;
wire uc_2023;
wire uc_2024;
wire uc_2025;
wire uc_2026;
wire uc_2027;
wire uc_2028;
wire uc_2029;
wire uc_2030;
wire uc_2031;
wire uc_2032;
wire uc_2033;
wire uc_2034;
wire uc_2035;
wire uc_2036;
wire uc_2037;
wire uc_2038;
wire uc_2039;
wire uc_2040;
wire uc_2041;
wire uc_2042;
wire uc_2043;
wire uc_2044;
wire uc_2045;
wire uc_2046;
wire uc_2047;
wire uc_2048;
wire uc_2049;
wire uc_2050;
wire uc_2051;
wire uc_2052;
wire uc_2053;
wire uc_2054;
wire uc_2055;
wire uc_2056;
wire uc_2057;
wire uc_2058;
wire uc_2059;
wire uc_2060;
wire uc_2061;
wire uc_2062;
wire uc_2063;
wire uc_2064;
wire uc_2065;
wire uc_2066;
wire uc_2067;
wire uc_2068;
wire uc_2069;
wire uc_2070;
wire uc_2071;
wire uc_2072;
wire uc_2073;
wire uc_2074;
wire uc_2075;
wire uc_2076;
wire uc_2077;
wire uc_2078;
wire uc_2079;
wire uc_2080;
wire uc_2081;
wire uc_2082;
wire uc_2083;
wire uc_2084;
wire uc_2085;
wire uc_2086;
wire uc_2087;
wire uc_2088;
wire uc_2089;
wire uc_2090;
wire uc_2091;
wire uc_2092;
wire uc_2093;
wire uc_2094;
wire uc_2095;
wire uc_2096;
wire uc_2097;
wire uc_2098;
wire uc_2099;
wire uc_2100;
wire uc_2101;
wire uc_2102;
wire uc_2103;
wire uc_2104;
wire uc_2105;
wire uc_2106;
wire uc_2107;
wire uc_2108;
wire uc_2109;
wire uc_2110;
wire uc_2111;
wire uc_2112;
wire uc_2113;
wire uc_2114;
wire uc_2115;
wire uc_2116;
wire uc_2117;
wire uc_2118;
wire uc_2119;
wire uc_2120;
wire uc_2121;
wire uc_2122;
wire uc_2123;
wire uc_2124;
wire uc_2125;
wire uc_2126;
wire uc_2127;
wire uc_2128;
wire uc_2129;
wire uc_2130;
wire uc_2131;
wire uc_2132;
wire uc_2133;
wire uc_2134;
wire uc_2135;
wire uc_2136;
wire uc_2137;
wire uc_2138;
wire uc_2139;
wire uc_2140;
wire uc_2141;
wire uc_2142;
wire uc_2143;
wire uc_2144;
wire uc_2145;
wire uc_2146;
wire uc_2147;
wire uc_2148;
wire uc_2149;
wire uc_2150;
wire uc_2151;
wire uc_2152;
wire uc_2153;
wire uc_2154;
wire uc_2155;
wire uc_2156;
wire uc_2157;
wire uc_2158;
wire uc_2159;
wire uc_2160;
wire uc_2161;
wire uc_2162;
wire uc_2163;
wire uc_2164;
wire uc_2165;
wire uc_2166;
wire uc_2167;
wire uc_2168;
wire uc_2169;
wire uc_2170;
wire uc_2171;
wire uc_2172;
wire uc_2173;
wire uc_2174;
wire uc_2175;
wire uc_2176;
wire uc_2177;
wire uc_2178;
wire uc_2179;
wire uc_2180;
wire uc_2181;
wire uc_2182;
wire uc_2183;
wire uc_2184;
wire uc_2185;
wire uc_2186;
wire uc_2187;
wire uc_2188;
wire uc_2189;
wire uc_2190;
wire uc_2191;
wire uc_2192;
wire uc_2193;
wire uc_2194;
wire uc_2195;
wire uc_2196;
wire uc_2197;
wire uc_2198;
wire uc_2199;
wire uc_2200;
wire uc_2201;
wire uc_2202;
wire uc_2203;
wire uc_2204;
wire uc_2205;
wire uc_2206;
wire uc_2207;
wire uc_2208;
wire uc_2209;
wire uc_2210;
wire uc_2211;
wire uc_2212;
wire uc_2213;
wire uc_2214;
wire uc_2215;
wire uc_2216;
wire uc_2217;
wire uc_2218;
wire uc_2219;
wire uc_2220;
wire uc_2221;
wire uc_2222;
wire uc_2223;
wire uc_2224;
wire uc_2225;
wire uc_2226;
wire uc_2227;
wire uc_2228;
wire uc_2229;
wire uc_2230;
wire uc_2231;
wire uc_2232;
wire uc_2233;
wire uc_2234;
wire uc_2235;
wire uc_2236;
wire uc_2237;
wire uc_2238;
wire uc_2239;
wire uc_2240;
wire uc_2241;
wire uc_2242;
wire uc_2243;
wire uc_2244;
wire uc_2245;
wire uc_2246;
wire uc_2247;
wire uc_2248;
wire uc_2249;
wire uc_2250;
wire uc_2251;
wire uc_2252;
wire uc_2253;
wire uc_2254;
wire uc_2255;
wire uc_2256;
wire uc_2257;
wire uc_2258;
wire uc_2259;
wire uc_2260;
wire uc_2261;
wire uc_2262;
wire uc_2263;
wire uc_2264;
wire uc_2265;
wire uc_2266;
wire uc_2267;
wire uc_2268;
wire uc_2269;
wire uc_2270;
wire uc_2271;
wire uc_2272;
wire uc_2273;
wire uc_2274;
wire uc_2275;
wire uc_2276;
wire uc_2277;
wire uc_2278;
wire uc_2279;
wire uc_2280;
wire uc_2281;
wire uc_2282;
wire uc_2283;
wire uc_2284;
wire uc_2285;
wire uc_2286;
wire uc_2287;
wire uc_2288;
wire uc_2289;
wire uc_2290;
wire uc_2291;
wire uc_2292;
wire uc_2293;
wire uc_2294;
wire uc_2295;
wire uc_2296;
wire uc_2297;
wire uc_2298;
wire uc_2299;
wire uc_2300;
wire uc_2301;
wire uc_2302;
wire uc_2303;
wire uc_2304;
wire uc_2305;
wire uc_2306;
wire uc_2307;
wire uc_2308;
wire uc_2309;
wire uc_2310;
wire uc_2311;
wire uc_2312;
wire uc_2313;
wire uc_2314;
wire uc_2315;
wire uc_2316;
wire uc_2317;
wire uc_2318;
wire uc_2319;
wire uc_2320;
wire uc_2321;
wire uc_2322;
wire uc_2323;
wire uc_2324;
wire uc_2325;
wire uc_2326;
wire uc_2327;
wire uc_2328;
wire uc_2329;
wire uc_2330;
wire uc_2331;
wire uc_2332;
wire uc_2333;
wire uc_2334;
wire uc_2335;
wire uc_2336;
wire uc_2337;
wire uc_2338;
wire uc_2339;
wire uc_2340;
wire uc_2341;
wire uc_2342;
wire uc_2343;
wire uc_2344;
wire uc_2345;
wire uc_2346;
wire uc_2347;
wire uc_2348;
wire uc_2349;
wire uc_2350;
wire uc_2351;
wire uc_2352;
wire uc_2353;
wire uc_2354;
wire uc_2355;
wire uc_2356;
wire uc_2357;
wire uc_2358;
wire uc_2359;
wire uc_2360;
wire uc_2361;
wire uc_2362;
wire uc_2363;
wire uc_2364;
wire uc_2365;
wire uc_2366;
wire uc_2367;
wire uc_2368;
wire uc_2369;
wire uc_2370;
wire uc_2371;
wire uc_2372;
wire uc_2373;
wire uc_2374;
wire uc_2375;
wire uc_2376;
wire uc_2377;
wire uc_2378;
wire uc_2379;
wire uc_2380;
wire uc_2381;
wire uc_2382;
wire uc_2383;
wire uc_2384;
wire uc_2385;
wire uc_2386;
wire uc_2387;
wire uc_2388;
wire uc_2389;
wire uc_2390;
wire uc_2391;
wire uc_2392;
wire uc_2393;
wire uc_2394;
wire uc_2395;
wire uc_2396;
wire uc_2397;
wire uc_2398;
wire uc_2399;
wire uc_2400;
wire uc_2401;
wire uc_2402;
wire uc_2403;
wire uc_2404;
wire uc_2405;
wire uc_2406;
wire uc_2407;
wire uc_2408;
wire uc_2409;
wire uc_2410;
wire uc_2411;
wire uc_2412;
wire uc_2413;
wire uc_2414;
wire uc_2415;
wire uc_2416;
wire uc_2417;
wire uc_2418;
wire uc_2419;
wire uc_2420;
wire uc_2421;
wire uc_2422;
wire uc_2423;
wire uc_2424;
wire uc_2425;
wire uc_2426;
wire uc_2427;
wire uc_2428;
wire uc_2429;
wire uc_2430;
wire uc_2431;
wire uc_2432;
wire uc_2433;
wire uc_2434;
wire uc_2435;
wire uc_2436;
wire uc_2437;
wire uc_2438;
wire uc_2439;
wire uc_2440;
wire uc_2441;
wire uc_2442;
wire uc_2443;
wire uc_2444;
wire uc_2445;
wire uc_2446;
wire uc_2447;
wire uc_2448;
wire uc_2449;
wire uc_2450;
wire uc_2451;
wire uc_2452;
wire uc_2453;
wire uc_2454;
wire uc_2455;
wire uc_2456;
wire uc_2457;
wire uc_2458;
wire uc_2459;
wire uc_2460;
wire uc_2461;
wire uc_2462;
wire uc_2463;
wire uc_2464;
wire uc_2465;
wire uc_2466;
wire uc_2467;
wire uc_2468;
wire uc_2469;
wire uc_2470;
wire uc_2471;
wire uc_2472;
wire uc_2473;
wire uc_2474;
wire uc_2475;
wire uc_2476;
wire uc_2477;
wire uc_2478;
wire uc_2479;
wire uc_2480;
wire uc_2481;
wire uc_2482;
wire uc_2483;
wire uc_2484;
wire uc_2485;
wire uc_2486;
wire uc_2487;
wire uc_2488;
wire uc_2489;
wire uc_2490;
wire uc_2491;
wire uc_2492;
wire uc_2493;
wire uc_2494;
wire uc_2495;
wire uc_2496;
wire uc_2497;
wire uc_2498;
wire uc_2499;
wire uc_2500;
wire uc_2501;
wire uc_2502;
wire uc_2503;
wire uc_2504;
wire uc_2505;
wire uc_2506;
wire uc_2507;
wire uc_2508;
wire uc_2509;
wire uc_2510;
wire uc_2511;
wire uc_2512;
wire uc_2513;
wire uc_2514;
wire uc_2515;
wire uc_2516;
wire uc_2517;
wire uc_2518;
wire uc_2519;
wire uc_2520;
wire uc_2521;
wire uc_2522;
wire uc_2523;
wire uc_2524;
wire uc_2525;
wire uc_2526;
wire uc_2527;
wire uc_2528;
wire uc_2529;
wire uc_2530;
wire uc_2531;
wire uc_2532;
wire uc_2533;
wire uc_2534;
wire uc_2535;
wire uc_2536;
wire uc_2537;
wire uc_2538;
wire uc_2539;
wire uc_2540;
wire uc_2541;
wire uc_2542;
wire uc_2543;
wire uc_2544;
wire uc_2545;
wire uc_2546;
wire uc_2547;
wire uc_2548;
wire uc_2549;
wire uc_2550;
wire uc_2551;
wire uc_2552;
wire uc_2553;
wire uc_2554;
wire uc_2555;
wire uc_2556;
wire uc_2557;
wire uc_2558;
wire uc_2559;
wire uc_2560;
wire uc_2561;
wire uc_2562;
wire uc_2563;
wire uc_2564;
wire uc_2565;
wire uc_2566;
wire uc_2567;
wire uc_2568;
wire uc_2569;
wire uc_2570;
wire uc_2571;
wire uc_2572;
wire uc_2573;
wire uc_2574;
wire uc_2575;
wire uc_2576;
wire uc_2577;
wire uc_2578;
wire uc_2579;
wire uc_2580;
wire uc_2581;
wire uc_2582;
wire uc_2583;
wire uc_2584;
wire uc_2585;
wire uc_2586;
wire uc_2587;
wire uc_2588;
wire uc_2589;
wire uc_2590;
wire uc_2591;
wire uc_2592;
wire uc_2593;
wire uc_2594;
wire uc_2595;
wire uc_2596;
wire uc_2597;
wire uc_2598;
wire uc_2599;
wire uc_2600;
wire uc_2601;
wire uc_2602;
wire uc_2603;
wire uc_2604;
wire uc_2605;
wire uc_2606;
wire uc_2607;
wire uc_2608;
wire uc_2609;
wire uc_2610;
wire uc_2611;
wire uc_2612;
wire uc_2613;
wire uc_2614;
wire uc_2615;
wire uc_2616;
wire uc_2617;
wire uc_2618;
wire uc_2619;
wire uc_2620;
wire uc_2621;
wire uc_2622;
wire uc_2623;
wire uc_2624;
wire uc_2625;
wire uc_2626;
wire uc_2627;
wire uc_2628;
wire uc_2629;
wire uc_2630;
wire uc_2631;
wire uc_2632;
wire uc_2633;
wire uc_2634;
wire uc_2635;
wire uc_2636;
wire uc_2637;
wire uc_2638;
wire uc_2639;
wire uc_2640;
wire uc_2641;
wire uc_2642;
wire uc_2643;
wire uc_2644;
wire uc_2645;
wire uc_2646;
wire uc_2647;
wire uc_2648;
wire uc_2649;
wire uc_2650;
wire uc_2651;
wire uc_2652;
wire uc_2653;
wire uc_2654;
wire uc_2655;
wire uc_2656;
wire uc_2657;
wire uc_2658;
wire uc_2659;
wire uc_2660;
wire uc_2661;
wire uc_2662;
wire uc_2663;
wire uc_2664;
wire uc_2665;
wire uc_2666;
wire uc_2667;
wire uc_2668;
wire uc_2669;
wire uc_2670;
wire uc_2671;
wire uc_2672;
wire uc_2673;
wire uc_2674;
wire uc_2675;
wire uc_2676;
wire uc_2677;
wire uc_2678;
wire uc_2679;
wire uc_2680;
wire uc_2681;
wire uc_2682;
wire uc_2683;
wire uc_2684;
wire uc_2685;
wire uc_2686;
wire uc_2687;
wire uc_2688;
wire uc_2689;
wire uc_2690;
wire uc_2691;
wire uc_2692;
wire uc_2693;
wire uc_2694;
wire uc_2695;
wire uc_2696;
wire uc_2697;
wire uc_2698;
wire uc_2699;
wire uc_2700;
wire uc_2701;
wire uc_2702;
wire uc_2703;
wire uc_2704;
wire uc_2705;
wire uc_2706;
wire uc_2707;
wire uc_2708;
wire uc_2709;
wire uc_2710;
wire uc_2711;
wire uc_2712;
wire uc_2713;
wire uc_2714;
wire uc_2715;
wire uc_2716;
wire uc_2717;
wire uc_2718;
wire uc_2719;
wire uc_2720;
wire uc_2721;
wire uc_2722;
wire uc_2723;
wire uc_2724;
wire uc_2725;
wire uc_2726;
wire uc_2727;
wire uc_2728;
wire uc_2729;
wire uc_2730;
wire uc_2731;
wire uc_2732;
wire uc_2733;
wire uc_2734;
wire uc_2735;
wire uc_2736;
wire uc_2737;
wire uc_2738;
wire uc_2739;
wire uc_2740;
wire uc_2741;
wire uc_2742;
wire uc_2743;
wire uc_2744;
wire uc_2745;
wire uc_2746;
wire uc_2747;
wire uc_2748;
wire uc_2749;
wire uc_2750;
wire uc_2751;
wire uc_2752;
wire uc_2753;
wire uc_2754;
wire uc_2755;
wire uc_2756;
wire uc_2757;
wire uc_2758;
wire uc_2759;
wire uc_2760;
wire uc_2761;
wire uc_2762;
wire uc_2763;
wire uc_2764;
wire uc_2765;
wire uc_2766;
wire uc_2767;
wire uc_2768;
wire uc_2769;
wire uc_2770;
wire uc_2771;
wire uc_2772;
wire uc_2773;
wire uc_2774;
wire uc_2775;
wire uc_2776;
wire uc_2777;
wire uc_2778;
wire uc_2779;
wire uc_2780;
wire uc_2781;
wire uc_2782;
wire uc_2783;
wire uc_2784;
wire uc_2785;
wire uc_2786;
wire uc_2787;
wire uc_2788;
wire uc_2789;
wire uc_2790;
wire uc_2791;
wire uc_2792;
wire uc_2793;
wire uc_2794;
wire uc_2795;
wire uc_2796;
wire uc_2797;
wire uc_2798;
wire uc_2799;
wire uc_2800;
wire uc_2801;
wire uc_2802;
wire uc_2803;
wire uc_2804;
wire uc_2805;
wire uc_2806;
wire uc_2807;
wire uc_2808;
wire uc_2809;
wire uc_2810;
wire uc_2811;
wire uc_2812;
wire uc_2813;
wire uc_2814;
wire uc_2815;
wire uc_2816;
wire uc_2817;
wire uc_2818;
wire uc_2819;
wire uc_2820;
wire uc_2821;
wire uc_2822;
wire uc_2823;
wire uc_2824;
wire uc_2825;
wire uc_2826;
wire uc_2827;
wire uc_2828;
wire uc_2829;
wire uc_2830;
wire uc_2831;
wire uc_2832;
wire uc_2833;
wire uc_2834;
wire uc_2835;
wire uc_2836;
wire uc_2837;
wire uc_2838;
wire uc_2839;
wire uc_2840;
wire uc_2841;
wire uc_2842;
wire uc_2843;
wire uc_2844;
wire uc_2845;
wire uc_2846;
wire uc_2847;
wire uc_2848;
wire uc_2849;
wire uc_2850;
wire uc_2851;
wire uc_2852;
wire uc_2853;
wire uc_2854;
wire uc_2855;
wire uc_2856;
wire uc_2857;
wire uc_2858;
wire uc_2859;
wire uc_2860;
wire uc_2861;
wire uc_2862;
wire uc_2863;
wire uc_2864;
wire uc_2865;
wire uc_2866;
wire uc_2867;
wire uc_2868;
wire uc_2869;
wire uc_2870;
wire uc_2871;
wire uc_2872;
wire uc_2873;
wire uc_2874;
wire uc_2875;
wire uc_2876;
wire uc_2877;
wire uc_2878;
wire uc_2879;
wire uc_2880;
wire uc_2881;
wire uc_2882;
wire uc_2883;
wire uc_2884;
wire uc_2885;
wire uc_2886;
wire uc_2887;
wire uc_2888;
wire uc_2889;
wire uc_2890;
wire uc_2891;
wire uc_2892;
wire uc_2893;
wire uc_2894;
wire uc_2895;
wire uc_2896;
wire uc_2897;
wire uc_2898;
wire uc_2899;
wire uc_2900;
wire uc_2901;
wire uc_2902;
wire uc_2903;
wire uc_2904;
wire uc_2905;
wire uc_2906;
wire uc_2907;
wire uc_2908;
wire uc_2909;
wire uc_2910;
wire uc_2911;
wire uc_2912;
wire uc_2913;
wire uc_2914;
wire uc_2915;
wire uc_2916;
wire uc_2917;
wire uc_2918;
wire uc_2919;
wire uc_2920;
wire uc_2921;
wire uc_2922;
wire uc_2923;
wire uc_2924;
wire uc_2925;
wire uc_2926;
wire uc_2927;
wire uc_2928;
wire uc_2929;
wire uc_2930;
wire uc_2931;
wire uc_2932;
wire uc_2933;
wire uc_2934;
wire uc_2935;
wire uc_2936;
wire uc_2937;
wire uc_2938;
wire uc_2939;
wire uc_2940;
wire uc_2941;
wire uc_2942;
wire uc_2943;
wire uc_2944;
wire uc_2945;
wire uc_2946;
wire uc_2947;
wire uc_2948;
wire uc_2949;
wire uc_2950;
wire uc_2951;
wire uc_2952;
wire uc_2953;
wire uc_2954;
wire uc_2955;
wire uc_2956;
wire uc_2957;
wire uc_2958;
wire uc_2959;
wire uc_2960;
wire uc_2961;
wire uc_2962;
wire uc_2963;
wire uc_2964;
wire uc_2965;
wire uc_2966;
wire uc_2967;
wire uc_2968;
wire uc_2969;
wire uc_2970;
wire uc_2971;
wire uc_2972;
wire uc_2973;
wire uc_2974;
wire uc_2975;
wire uc_2976;
wire uc_2977;
wire uc_2978;
wire uc_2979;
wire uc_2980;
wire uc_2981;
wire uc_2982;
wire uc_2983;
wire uc_2984;
wire uc_2985;
wire uc_2986;
wire uc_2987;
wire uc_2988;
wire uc_2989;
wire uc_2990;
wire uc_2991;
wire uc_2992;
wire uc_2993;
wire uc_2994;
wire uc_2995;
wire uc_2996;
wire uc_2997;
wire uc_2998;
wire uc_2999;
wire uc_3000;
wire uc_3001;
wire uc_3002;
wire uc_3003;
wire uc_3004;
wire uc_3005;
wire uc_3006;
wire uc_3007;
wire uc_3008;
wire uc_3009;
wire uc_3010;
wire uc_3011;
wire uc_3012;
wire uc_3013;
wire uc_3014;
wire uc_3015;
wire uc_3016;
wire uc_3017;
wire uc_3018;
wire uc_3019;
wire uc_3020;
wire uc_3021;
wire uc_3022;
wire uc_3023;
wire uc_3024;
wire uc_3025;
wire uc_3026;
wire uc_3027;
wire uc_3028;
wire uc_3029;
wire uc_3030;
wire uc_3031;
wire uc_3032;
wire uc_3033;
wire uc_3034;
wire uc_3035;
wire uc_3036;
wire uc_3037;
wire uc_3038;
wire uc_3039;
wire uc_3040;
wire uc_3041;
wire uc_3042;
wire uc_3043;
wire uc_3044;
wire uc_3045;
wire uc_3046;
wire uc_3047;
wire uc_3048;
wire uc_3049;
wire uc_3050;
wire uc_3051;
wire uc_3052;
wire uc_3053;
wire uc_3054;
wire uc_3055;
wire uc_3056;
wire uc_3057;
wire uc_3058;
wire uc_3059;
wire uc_3060;
wire uc_3061;
wire uc_3062;
wire uc_3063;
wire uc_3064;
wire uc_3065;
wire uc_3066;
wire uc_3067;
wire uc_3068;
wire uc_3069;
wire uc_3070;
wire uc_3071;
wire uc_3072;
wire uc_3073;
wire uc_3074;
wire uc_3075;
wire uc_3076;
wire uc_3077;
wire uc_3078;
wire uc_3079;
wire uc_3080;
wire uc_3081;
wire uc_3082;
wire uc_3083;
wire uc_3084;
wire uc_3085;
wire uc_3086;
wire uc_3087;
wire uc_3088;
wire uc_3089;
wire uc_3090;
wire uc_3091;
wire uc_3092;
wire uc_3093;
wire uc_3094;
wire uc_3095;
wire uc_3096;
wire uc_3097;
wire uc_3098;
wire uc_3099;
wire uc_3100;
wire uc_3101;
wire uc_3102;
wire uc_3103;
wire uc_3104;
wire uc_3105;
wire uc_3106;
wire uc_3107;
wire uc_3108;
wire uc_3109;
wire uc_3110;
wire uc_3111;
wire uc_3112;
wire uc_3113;
wire uc_3114;
wire uc_3115;
wire uc_3116;
wire uc_3117;
wire uc_3118;
wire uc_3119;
wire uc_3120;
wire uc_3121;
wire uc_3122;
wire uc_3123;
wire uc_3124;
wire uc_3125;
wire uc_3126;
wire uc_3127;
wire uc_3128;
wire uc_3129;
wire uc_3130;
wire uc_3131;
wire uc_3132;
wire uc_3133;
wire uc_3134;
wire uc_3135;
wire uc_3136;
wire uc_3137;
wire uc_3138;
wire uc_3139;
wire uc_3140;
wire uc_3141;
wire uc_3142;
wire uc_3143;
wire uc_3144;
wire uc_3145;
wire uc_3146;
wire uc_3147;
wire uc_3148;
wire uc_3149;
wire uc_3150;
wire uc_3151;
wire uc_3152;
wire uc_3153;
wire uc_3154;
wire uc_3155;
wire uc_3156;
wire uc_3157;
wire uc_3158;
wire uc_3159;
wire uc_3160;
wire uc_3161;
wire uc_3162;
wire uc_3163;
wire uc_3164;
wire uc_3165;
wire uc_3166;
wire uc_3167;
wire uc_3168;
wire uc_3169;
wire uc_3170;
wire uc_3171;
wire uc_3172;
wire uc_3173;
wire uc_3174;
wire uc_3175;
wire uc_3176;
wire uc_3177;
wire uc_3178;
wire uc_3179;
wire uc_3180;
wire uc_3181;
wire uc_3182;
wire uc_3183;
wire uc_3184;
wire uc_3185;
wire uc_3186;
wire uc_3187;
wire uc_3188;
wire uc_3189;
wire uc_3190;
wire uc_3191;
wire uc_3192;
wire uc_3193;
wire uc_3194;
wire uc_3195;
wire uc_3196;
wire uc_3197;
wire uc_3198;
wire uc_3199;
wire uc_3200;
wire uc_3201;
wire uc_3202;
wire uc_3203;
wire uc_3204;
wire uc_3205;
wire uc_3206;
wire uc_3207;
wire uc_3208;
wire uc_3209;
wire uc_3210;
wire uc_3211;
wire uc_3212;
wire uc_3213;
wire uc_3214;
wire uc_3215;
wire uc_3216;
wire uc_3217;
wire uc_3218;
wire uc_3219;
wire uc_3220;
wire uc_3221;
wire uc_3222;
wire uc_3223;
wire uc_3224;
wire uc_3225;
wire uc_3226;
wire uc_3227;
wire uc_3228;
wire uc_3229;
wire uc_3230;
wire uc_3231;
wire uc_3232;
wire uc_3233;
wire uc_3234;
wire uc_3235;
wire uc_3236;
wire uc_3237;
wire uc_3238;
wire uc_3239;
wire uc_3240;
wire uc_3241;
wire uc_3242;
wire uc_3243;
wire uc_3244;
wire uc_3245;
wire uc_3246;
wire uc_3247;
wire uc_3248;
wire uc_3249;
wire uc_3250;
wire uc_3251;
wire uc_3252;
wire uc_3253;
wire uc_3254;
wire uc_3255;
wire uc_3256;
wire uc_3257;
wire uc_3258;
wire uc_3259;
wire uc_3260;
wire uc_3261;
wire uc_3262;
wire uc_3263;
wire uc_3264;
wire uc_3265;
wire uc_3266;
wire uc_3267;
wire uc_3268;
wire uc_3269;
wire uc_3270;
wire uc_3271;
wire uc_3272;
wire uc_3273;
wire uc_3274;
wire uc_3275;
wire uc_3276;
wire uc_3277;
wire uc_3278;
wire uc_3279;
wire uc_3280;
wire uc_3281;
wire uc_3282;
wire uc_3283;
wire uc_3284;
wire uc_3285;
wire uc_3286;
wire uc_3287;
wire uc_3288;
wire uc_3289;
wire uc_3290;
wire uc_3291;
wire uc_3292;
wire uc_3293;
wire uc_3294;
wire uc_3295;
wire uc_3296;
wire uc_3297;
wire uc_3298;
wire uc_3299;
wire uc_3300;
wire uc_3301;
wire uc_3302;
wire uc_3303;
wire uc_3304;
wire uc_3305;
wire uc_3306;
wire uc_3307;
wire uc_3308;
wire uc_3309;
wire uc_3310;
wire uc_3311;
wire uc_3312;
wire uc_3313;
wire uc_3314;
wire uc_3315;
wire uc_3316;
wire uc_3317;
wire uc_3318;
wire uc_3319;
wire uc_3320;
wire uc_3321;
wire uc_3322;
wire uc_3323;
wire uc_3324;
wire uc_3325;
wire uc_3326;
wire uc_3327;
wire uc_3328;
wire uc_3329;
wire uc_3330;
wire uc_3331;
wire uc_3332;
wire uc_3333;
wire uc_3334;
wire uc_3335;
wire uc_3336;
wire uc_3337;
wire uc_3338;
wire uc_3339;
wire uc_3340;
wire uc_3341;
wire uc_3342;
wire uc_3343;
wire uc_3344;
wire uc_3345;
wire uc_3346;
wire uc_3347;
wire uc_3348;
wire uc_3349;
wire uc_3350;
wire uc_3351;
wire uc_3352;
wire uc_3353;
wire uc_3354;
wire uc_3355;
wire uc_3356;
wire uc_3357;
wire uc_3358;
wire uc_3359;
wire uc_3360;
wire uc_3361;
wire uc_3362;
wire uc_3363;
wire uc_3364;
wire uc_3365;
wire uc_3366;
wire uc_3367;
wire uc_3368;
wire uc_3369;
wire uc_3370;
wire uc_3371;
wire uc_3372;
wire uc_3373;
wire uc_3374;
wire uc_3375;
wire uc_3376;
wire uc_3377;
wire uc_3378;
wire uc_3379;
wire uc_3380;
wire uc_3381;
wire uc_3382;
wire uc_3383;
wire uc_3384;
wire uc_3385;
wire uc_3386;
wire uc_3387;
wire uc_3388;
wire uc_3389;
wire uc_3390;
wire uc_3391;
wire uc_3392;
wire uc_3393;
wire uc_3394;
wire uc_3395;
wire uc_3396;
wire uc_3397;
wire uc_3398;
wire uc_3399;
wire uc_3400;
wire uc_3401;
wire uc_3402;
wire uc_3403;
wire uc_3404;
wire uc_3405;
wire uc_3406;
wire uc_3407;
wire uc_3408;
wire uc_3409;
wire uc_3410;
wire uc_3411;
wire uc_3412;
wire uc_3413;
wire uc_3414;
wire uc_3415;
wire uc_3416;
wire uc_3417;
wire uc_3418;
wire uc_3419;
wire uc_3420;
wire uc_3421;
wire uc_3422;
wire uc_3423;
wire uc_3424;
wire uc_3425;
wire uc_3426;
wire uc_3427;
wire uc_3428;
wire uc_3429;
wire uc_3430;
wire uc_3431;
wire uc_3432;
wire uc_3433;
wire uc_3434;
wire uc_3435;
wire uc_3436;
wire uc_3437;
wire uc_3438;
wire uc_3439;
wire uc_3440;
wire uc_3441;
wire uc_3442;
wire uc_3443;
wire uc_3444;
wire uc_3445;
wire uc_3446;
wire uc_3447;
wire uc_3448;
wire uc_3449;
wire uc_3450;
wire uc_3451;
wire uc_3452;
wire uc_3453;
wire uc_3454;
wire uc_3455;
wire uc_3456;
wire uc_3457;
wire uc_3458;
wire uc_3459;
wire uc_3460;
wire uc_3461;
wire uc_3462;
wire uc_3463;
wire uc_3464;
wire uc_3465;
wire uc_3466;
wire uc_3467;
wire uc_3468;
wire uc_3469;
wire uc_3470;
wire uc_3471;
wire uc_3472;
wire uc_3473;
wire uc_3474;
wire uc_3475;
wire uc_3476;
wire uc_3477;
wire uc_3478;
wire uc_3479;
wire uc_3480;
wire uc_3481;
wire uc_3482;
wire uc_3483;
wire uc_3484;
wire uc_3485;
wire uc_3486;
wire uc_3487;
wire uc_3488;
wire uc_3489;
wire uc_3490;
wire uc_3491;
wire uc_3492;
wire uc_3493;
wire uc_3494;
wire uc_3495;
wire uc_3496;
wire uc_3497;
wire uc_3498;
wire uc_3499;
wire uc_3500;
wire uc_3501;
wire uc_3502;
wire uc_3503;
wire uc_3504;
wire uc_3505;
wire uc_3506;
wire uc_3507;
wire uc_3508;
wire uc_3509;
wire uc_3510;
wire uc_3511;
wire uc_3512;
wire uc_3513;
wire uc_3514;
wire uc_3515;
wire uc_3516;
wire uc_3517;
wire uc_3518;
wire uc_3519;
wire uc_3520;
wire uc_3521;
wire uc_3522;
wire uc_3523;
wire uc_3524;
wire uc_3525;
wire uc_3526;
wire uc_3527;
wire uc_3528;
wire uc_3529;
wire uc_3530;
wire uc_3531;
wire uc_3532;
wire uc_3533;
wire uc_3534;
wire uc_3535;
wire uc_3536;
wire uc_3537;
wire uc_3538;
wire uc_3539;
wire uc_3540;
wire uc_3541;
wire uc_3542;
wire uc_3543;
wire uc_3544;
wire uc_3545;
wire uc_3546;
wire uc_3547;
wire uc_3548;
wire uc_3549;
wire uc_3550;
wire uc_3551;
wire uc_3552;
wire uc_3553;
wire uc_3554;
wire uc_3555;
wire uc_3556;
wire uc_3557;
wire uc_3558;
wire uc_3559;
wire uc_3560;
wire uc_3561;
wire uc_3562;
wire uc_3563;
wire uc_3564;
wire uc_3565;
wire uc_3566;
wire uc_3567;
wire uc_3568;
wire uc_3569;
wire uc_3570;
wire uc_3571;
wire uc_3572;
wire uc_3573;
wire uc_3574;
wire uc_3575;
wire uc_3576;
wire uc_3577;
wire uc_3578;
wire uc_3579;
wire uc_3580;
wire uc_3581;
wire uc_3582;
wire uc_3583;
wire uc_3584;
wire uc_3585;
wire uc_3586;
wire uc_3587;
wire uc_3588;
wire uc_3589;
wire uc_3590;
wire uc_3591;
wire uc_3592;
wire uc_3593;
wire uc_3594;
wire uc_3595;
wire uc_3596;
wire uc_3597;
wire uc_3598;
wire uc_3599;
wire uc_3600;
wire uc_3601;
wire uc_3602;
wire uc_3603;
wire uc_3604;
wire uc_3605;
wire uc_3606;
wire uc_3607;
wire uc_3608;
wire uc_3609;
wire uc_3610;
wire uc_3611;
wire uc_3612;
wire uc_3613;
wire uc_3614;
wire uc_3615;
wire uc_3616;
wire uc_3617;
wire uc_3618;
wire uc_3619;
wire uc_3620;
wire uc_3621;
wire uc_3622;
wire uc_3623;
wire uc_3624;
wire uc_3625;
wire uc_3626;
wire uc_3627;
wire uc_3628;
wire uc_3629;
wire uc_3630;
wire uc_3631;
wire uc_3632;
wire uc_3633;
wire uc_3634;
wire uc_3635;
wire uc_3636;
wire uc_3637;
wire uc_3638;
wire uc_3639;
wire uc_3640;
wire uc_3641;
wire uc_3642;
wire uc_3643;
wire uc_3644;
wire uc_3645;
wire uc_3646;
wire uc_3647;
wire uc_3648;
wire uc_3649;
wire uc_3650;
wire uc_3651;
wire uc_3652;
wire uc_3653;
wire uc_3654;
wire uc_3655;
wire uc_3656;
wire uc_3657;
wire uc_3658;
wire uc_3659;
wire uc_3660;
wire uc_3661;
wire uc_3662;
wire uc_3663;
wire uc_3664;
wire uc_3665;
wire uc_3666;
wire uc_3667;
wire uc_3668;
wire uc_3669;
wire uc_3670;
wire uc_3671;
wire uc_3672;
wire uc_3673;
wire uc_3674;
wire uc_3675;
wire uc_3676;
wire uc_3677;
wire uc_3678;
wire uc_3679;
wire uc_3680;
wire uc_3681;
wire uc_3682;
wire uc_3683;
wire uc_3684;
wire uc_3685;
wire uc_3686;
wire uc_3687;
wire uc_3688;
wire uc_3689;
wire uc_3690;
wire uc_3691;
wire uc_3692;
wire uc_3693;
wire uc_3694;
wire uc_3695;
wire uc_3696;
wire uc_3697;
wire uc_3698;
wire uc_3699;
wire uc_3700;
wire uc_3701;
wire uc_3702;
wire uc_3703;
wire uc_3704;
wire uc_3705;
wire uc_3706;
wire uc_3707;
wire uc_3708;
wire uc_3709;
wire uc_3710;
wire uc_3711;
wire uc_3712;
wire uc_3713;
wire uc_3714;
wire uc_3715;
wire uc_3716;
wire uc_3717;
wire uc_3718;
wire uc_3719;
wire uc_3720;
wire uc_3721;
wire uc_3722;
wire uc_3723;
wire uc_3724;
wire uc_3725;
wire uc_3726;
wire uc_3727;
wire uc_3728;
wire uc_3729;
wire uc_3730;
wire uc_3731;
wire uc_3732;
wire uc_3733;
wire uc_3734;
wire uc_3735;
wire uc_3736;
wire uc_3737;
wire uc_3738;
wire uc_3739;
wire uc_3740;
wire uc_3741;
wire uc_3742;
wire uc_3743;
wire uc_3744;
wire uc_3745;
wire uc_3746;
wire uc_3747;
wire uc_3748;
wire uc_3749;
wire uc_3750;
wire uc_3751;
wire uc_3752;
wire uc_3753;
wire uc_3754;
wire uc_3755;
wire uc_3756;
wire uc_3757;
wire uc_3758;
wire uc_3759;
wire uc_3760;
wire uc_3761;
wire uc_3762;
wire uc_3763;
wire uc_3764;
wire uc_3765;
wire uc_3766;
wire uc_3767;
wire uc_3768;
wire uc_3769;
wire uc_3770;
wire uc_3771;
wire uc_3772;
wire uc_3773;
wire uc_3774;
wire uc_3775;
wire uc_3776;
wire uc_3777;
wire uc_3778;
wire uc_3779;
wire uc_3780;
wire uc_3781;
wire uc_3782;
wire uc_3783;
wire uc_3784;
wire uc_3785;
wire uc_3786;
wire uc_3787;
wire uc_3788;
wire uc_3789;
wire uc_3790;
wire uc_3791;
wire uc_3792;
wire uc_3793;
wire uc_3794;
wire uc_3795;
wire uc_3796;
wire uc_3797;
wire uc_3798;
wire uc_3799;
wire uc_3800;
wire uc_3801;
wire uc_3802;
wire uc_3803;
wire uc_3804;
wire uc_3805;
wire uc_3806;
wire uc_3807;
wire uc_3808;
wire uc_3809;
wire uc_3810;
wire uc_3811;
wire uc_3812;
wire uc_3813;
wire uc_3814;
wire uc_3815;
wire uc_3816;
wire uc_3817;
wire uc_3818;
wire uc_3819;
wire uc_3820;
wire uc_3821;
wire uc_3822;
wire uc_3823;
wire uc_3824;
wire uc_3825;
wire uc_3826;
wire uc_3827;
wire uc_3828;
wire uc_3829;
wire uc_3830;
wire uc_3831;
wire uc_3832;
wire uc_3833;
wire uc_3834;
wire uc_3835;
wire uc_3836;
wire uc_3837;
wire uc_3838;
wire uc_3839;
wire uc_3840;
wire uc_3841;
wire uc_3842;
wire uc_3843;
wire uc_3844;
wire uc_3845;
wire uc_3846;
wire uc_3847;
wire uc_3848;
wire uc_3849;
wire uc_3850;
wire uc_3851;
wire uc_3852;
wire uc_3853;
wire uc_3854;
wire uc_3855;
wire uc_3856;
wire uc_3857;
wire uc_3858;
wire uc_3859;
wire uc_3860;
wire uc_3861;
wire uc_3862;
wire uc_3863;
wire uc_3864;
wire uc_3865;
wire uc_3866;
wire uc_3867;
wire uc_3868;
wire uc_3869;
wire uc_3870;
wire uc_3871;
wire uc_3872;
wire uc_3873;
wire uc_3874;
wire uc_3875;
wire uc_3876;
wire uc_3877;
wire uc_3878;
wire uc_3879;
wire uc_3880;
wire uc_3881;
wire uc_3882;
wire uc_3883;
wire uc_3884;
wire uc_3885;
wire uc_3886;
wire uc_3887;
wire uc_3888;
wire uc_3889;
wire uc_3890;
wire uc_3891;
wire uc_3892;
wire uc_3893;
wire uc_3894;
wire uc_3895;
wire uc_3896;
wire uc_3897;
wire uc_3898;
wire uc_3899;
wire uc_3900;
wire uc_3901;
wire uc_3902;
wire uc_3903;
wire uc_3904;
wire uc_3905;
wire uc_3906;
wire uc_3907;
wire uc_3908;
wire uc_3909;
wire uc_3910;
wire uc_3911;
wire uc_3912;
wire uc_3913;
wire uc_3914;
wire uc_3915;
wire uc_3916;
wire uc_3917;
wire uc_3918;
wire uc_3919;
wire uc_3920;
wire uc_3921;
wire uc_3922;
wire uc_3923;
wire uc_3924;
wire uc_3925;
wire uc_3926;
wire uc_3927;
wire uc_3928;
wire uc_3929;
wire uc_3930;
wire uc_3931;
wire uc_3932;
wire uc_3933;
wire uc_3934;
wire uc_3935;
wire uc_3936;
wire uc_3937;
wire uc_3938;
wire uc_3939;
wire uc_3940;
wire uc_3941;
wire uc_3942;
wire uc_3943;
wire uc_3944;
wire uc_3945;
wire uc_3946;
wire uc_3947;
wire uc_3948;
wire uc_3949;
wire uc_3950;
wire uc_3951;
wire uc_3952;
wire uc_3953;
wire uc_3954;
wire uc_3955;
wire uc_3956;
wire uc_3957;
wire uc_3958;
wire uc_3959;
wire uc_3960;
wire uc_3961;
wire uc_3962;
wire uc_3963;
wire uc_3964;
wire uc_3965;
wire uc_3966;
wire uc_3967;
wire uc_3968;
wire uc_3969;
wire uc_3970;
wire uc_3971;
wire uc_3972;
wire uc_3973;
wire uc_3974;
wire uc_3975;
wire uc_3976;
wire uc_3977;
wire uc_3978;
wire uc_3979;
wire uc_3980;
wire uc_3981;
wire uc_3982;
wire uc_3983;
wire uc_3984;
wire uc_3985;
wire uc_3986;
wire uc_3987;
wire uc_3988;
wire uc_3989;
wire uc_3990;
wire uc_3991;
wire uc_3992;
wire uc_3993;
wire uc_3994;
wire uc_3995;
wire uc_3996;
wire uc_3997;
wire uc_3998;
wire uc_3999;
wire uc_4000;
wire uc_4001;
wire uc_4002;
wire uc_4003;
wire uc_4004;
wire uc_4005;
wire uc_4006;
wire uc_4007;
wire uc_4008;
wire uc_4009;
wire uc_4010;
wire uc_4011;
wire uc_4012;
wire uc_4013;
wire uc_4014;
wire uc_4015;
wire uc_4016;
wire uc_4017;
wire uc_4018;
wire uc_4019;
wire uc_4020;
wire uc_4021;
wire uc_4022;
wire uc_4023;
wire uc_4024;
wire uc_4025;
wire uc_4026;
wire uc_4027;
wire uc_4028;
wire uc_4029;
wire uc_4030;
wire uc_4031;
wire uc_4032;
wire uc_4033;
wire uc_4034;
wire uc_4035;
wire uc_4036;
wire uc_4037;
wire uc_4038;
wire uc_4039;
wire uc_4040;
wire uc_4041;
wire uc_4042;
wire uc_4043;
wire uc_4044;
wire uc_4045;
wire uc_4046;
wire uc_4047;
wire uc_4048;
wire uc_4049;
wire uc_4050;
wire uc_4051;
wire uc_4052;
wire uc_4053;
wire uc_4054;
wire uc_4055;
wire uc_4056;
wire uc_4057;
wire uc_4058;
wire uc_4059;
wire uc_4060;
wire uc_4061;
wire uc_4062;
wire uc_4063;
wire uc_4064;
wire uc_4065;
wire uc_4066;
wire uc_4067;
wire uc_4068;
wire uc_4069;
wire uc_4070;
wire uc_4071;
wire uc_4072;
wire uc_4073;
wire uc_4074;
wire uc_4075;
wire uc_4076;
wire uc_4077;
wire uc_4078;
wire uc_4079;
wire uc_4080;
wire uc_4081;
wire uc_4082;
wire uc_4083;
wire uc_4084;
wire uc_4085;
wire uc_4086;
wire uc_4087;
wire uc_4088;
wire uc_4089;
wire uc_4090;
wire uc_4091;
wire uc_4092;
wire uc_4093;
wire uc_4094;
wire uc_4095;
wire uc_4096;
wire uc_4097;
wire uc_4098;
wire uc_4099;
wire uc_4100;
wire uc_4101;
wire uc_4102;
wire uc_4103;
wire uc_4104;
wire uc_4105;
wire uc_4106;
wire uc_4107;
wire uc_4108;
wire uc_4109;
wire uc_4110;
wire uc_4111;
wire uc_4112;
wire uc_4113;
wire uc_4114;
wire uc_4115;
wire uc_4116;
wire uc_4117;
wire uc_4118;
wire uc_4119;
wire uc_4120;
wire uc_4121;
wire uc_4122;
wire uc_4123;
wire uc_4124;
wire uc_4125;
wire uc_4126;
wire uc_4127;
wire uc_4128;
wire uc_4129;
wire uc_4130;
wire uc_4131;
wire uc_4132;
wire uc_4133;
wire uc_4134;
wire uc_4135;
wire uc_4136;
wire uc_4137;
wire uc_4138;
wire uc_4139;
wire uc_4140;
wire uc_4141;
wire uc_4142;
wire uc_4143;
wire uc_4144;
wire uc_4145;
wire uc_4146;
wire uc_4147;
wire uc_4148;
wire uc_4149;
wire uc_4150;
wire uc_4151;
wire uc_4152;
wire uc_4153;
wire uc_4154;
wire uc_4155;
wire uc_4156;
wire uc_4157;
wire uc_4158;
wire uc_4159;
wire uc_4160;
wire uc_4161;
wire uc_4162;
wire uc_4163;
wire uc_4164;
wire uc_4165;
wire uc_4166;
wire uc_4167;
wire uc_4168;
wire uc_4169;
wire uc_4170;
wire uc_4171;
wire uc_4172;
wire uc_4173;
wire uc_4174;
wire uc_4175;
wire uc_4176;
wire uc_4177;
wire uc_4178;
wire uc_4179;
wire uc_4180;
wire uc_4181;
wire uc_4182;
wire uc_4183;
wire uc_4184;
wire uc_4185;
wire uc_4186;
wire uc_4187;
wire uc_4188;
wire uc_4189;
wire uc_4190;
wire uc_4191;
wire uc_4192;
wire uc_4193;
wire uc_4194;
wire uc_4195;
wire uc_4196;
wire uc_4197;
wire uc_4198;
wire uc_4199;
wire uc_4200;
wire uc_4201;
wire uc_4202;
wire uc_4203;
wire uc_4204;
wire uc_4205;
wire uc_4206;
wire uc_4207;
wire uc_4208;
wire uc_4209;
wire uc_4210;
wire uc_4211;
wire uc_4212;
wire uc_4213;
wire uc_4214;
wire uc_4215;
wire uc_4216;
wire uc_4217;
wire uc_4218;
wire uc_4219;
wire uc_4220;
wire uc_4221;
wire uc_4222;
wire uc_4223;
wire uc_4224;
wire uc_4225;
wire uc_4226;
wire uc_4227;
wire uc_4228;
wire uc_4229;
wire uc_4230;
wire uc_4231;
wire uc_4232;
wire uc_4233;
wire uc_4234;
wire uc_4235;
wire uc_4236;
wire uc_4237;
wire uc_4238;
wire uc_4239;
wire uc_4240;
wire uc_4241;
wire uc_4242;
wire uc_4243;
wire uc_4244;
wire uc_4245;
wire uc_4246;
wire uc_4247;
wire uc_4248;
wire uc_4249;
wire uc_4250;
wire uc_4251;
wire uc_4252;
wire uc_4253;
wire uc_4254;
wire uc_4255;
wire uc_4256;
wire uc_4257;
wire uc_4258;
wire uc_4259;
wire uc_4260;
wire uc_4261;
wire uc_4262;
wire uc_4263;
wire uc_4264;
wire uc_4265;
wire uc_4266;
wire uc_4267;
wire uc_4268;
wire uc_4269;
wire uc_4270;
wire uc_4271;
wire uc_4272;
wire uc_4273;
wire uc_4274;
wire uc_4275;
wire uc_4276;
wire uc_4277;
wire uc_4278;
wire uc_4279;
wire uc_4280;
wire uc_4281;
wire uc_4282;
wire uc_4283;
wire uc_4284;
wire uc_4285;
wire uc_4286;
wire uc_4287;
wire uc_4288;
wire uc_4289;
wire uc_4290;
wire uc_4291;
wire uc_4292;
wire uc_4293;
wire uc_4294;
wire uc_4295;
wire uc_4296;
wire uc_4297;
wire uc_4298;
wire uc_4299;
wire uc_4300;
wire uc_4301;
wire uc_4302;
wire uc_4303;
wire uc_4304;
wire uc_4305;
wire uc_4306;
wire uc_4307;
wire uc_4308;
wire uc_4309;
wire uc_4310;
wire uc_4311;
wire uc_4312;
wire uc_4313;
wire uc_4314;
wire uc_4315;
wire uc_4316;
wire uc_4317;
wire uc_4318;
wire uc_4319;
wire uc_4320;
wire uc_4321;
wire uc_4322;
wire uc_4323;
wire uc_4324;
wire uc_4325;
wire uc_4326;
wire uc_4327;
wire uc_4328;
wire uc_4329;
wire uc_4330;
wire uc_4331;
wire uc_4332;
wire uc_4333;
wire uc_4334;
wire uc_4335;
wire uc_4336;
wire uc_4337;
wire uc_4338;
wire uc_4339;
wire uc_4340;
wire uc_4341;
wire uc_4342;
wire uc_4343;
wire uc_4344;
wire uc_4345;
wire uc_4346;
wire uc_4347;
wire uc_4348;
wire uc_4349;
wire uc_4350;
wire uc_4351;
wire uc_4352;
wire uc_4353;
wire uc_4354;
wire uc_4355;
wire uc_4356;
wire uc_4357;
wire uc_4358;
wire uc_4359;
wire uc_4360;
wire uc_4361;
wire uc_4362;
wire uc_4363;
wire uc_4364;
wire uc_4365;
wire uc_4366;
wire uc_4367;
wire uc_4368;
wire uc_4369;
wire uc_4370;
wire uc_4371;
wire uc_4372;
wire uc_4373;
wire uc_4374;
wire uc_4375;
wire uc_4376;
wire uc_4377;
wire uc_4378;
wire uc_4379;
wire uc_4380;
wire uc_4381;
wire uc_4382;
wire uc_4383;
wire uc_4384;
wire uc_4385;
wire uc_4386;
wire uc_4387;
wire uc_4388;
wire uc_4389;
wire uc_4390;
wire uc_4391;
wire uc_4392;
wire uc_4393;
wire uc_4394;
wire uc_4395;
wire uc_4396;
wire uc_4397;
wire uc_4398;
wire uc_4399;
wire uc_4400;
wire uc_4401;
wire uc_4402;
wire uc_4403;
wire uc_4404;
wire uc_4405;
wire uc_4406;
wire uc_4407;
wire uc_4408;
wire uc_4409;
wire uc_4410;
wire uc_4411;
wire uc_4412;
wire uc_4413;
wire uc_4414;
wire uc_4415;
wire uc_4416;
wire uc_4417;
wire uc_4418;
wire uc_4419;
wire uc_4420;
wire uc_4421;
wire uc_4422;
wire uc_4423;
wire uc_4424;
wire uc_4425;
wire uc_4426;
wire uc_4427;
wire uc_4428;
wire uc_4429;
wire uc_4430;
wire uc_4431;
wire uc_4432;
wire uc_4433;
wire uc_4434;
wire uc_4435;
wire uc_4436;
wire uc_4437;
wire uc_4438;
wire uc_4439;
wire uc_4440;
wire uc_4441;
wire uc_4442;
wire uc_4443;
wire uc_4444;
wire uc_4445;
wire uc_4446;
wire uc_4447;
wire uc_4448;
wire uc_4449;
wire uc_4450;
wire uc_4451;
wire uc_4452;
wire uc_4453;
wire uc_4454;
wire uc_4455;
wire uc_4456;
wire uc_4457;
wire uc_4458;
wire uc_4459;
wire uc_4460;
wire uc_4461;
wire uc_4462;
wire uc_4463;
wire uc_4464;
wire uc_4465;
wire uc_4466;
wire uc_4467;
wire uc_4468;
wire uc_4469;
wire uc_4470;
wire uc_4471;
wire uc_4472;
wire uc_4473;
wire uc_4474;
wire uc_4475;
wire uc_4476;
wire uc_4477;
wire uc_4478;
wire uc_4479;
wire uc_4480;
wire uc_4481;
wire uc_4482;
wire uc_4483;
wire uc_4484;
wire uc_4485;
wire uc_4486;
wire uc_4487;
wire uc_4488;
wire uc_4489;
wire uc_4490;
wire uc_4491;
wire uc_4492;
wire uc_4493;
wire uc_4494;
wire uc_4495;
wire uc_4496;
wire uc_4497;
wire uc_4498;
wire uc_4499;
wire uc_4500;
wire uc_4501;
wire uc_4502;
wire uc_4503;
wire uc_4504;
wire uc_4505;
wire uc_4506;
wire uc_4507;
wire uc_4508;
wire uc_4509;
wire uc_4510;
wire uc_4511;
wire uc_4512;
wire uc_4513;
wire uc_4514;
wire uc_4515;
wire uc_4516;
wire uc_4517;
wire uc_4518;
wire uc_4519;
wire uc_4520;
wire uc_4521;
wire uc_4522;
wire uc_4523;
wire uc_4524;
wire uc_4525;
wire uc_4526;
wire uc_4527;
wire uc_4528;
wire uc_4529;
wire uc_4530;
wire uc_4531;
wire uc_4532;
wire uc_4533;
wire uc_4534;
wire uc_4535;
wire uc_4536;
wire uc_4537;
wire uc_4538;
wire uc_4539;
wire uc_4540;
wire uc_4541;
wire uc_4542;
wire uc_4543;
wire uc_4544;
wire uc_4545;
wire uc_4546;
wire uc_4547;
wire uc_4548;
wire uc_4549;
wire uc_4550;
wire uc_4551;
wire uc_4552;
wire uc_4553;
wire uc_4554;
wire uc_4555;
wire uc_4556;
wire uc_4557;
wire uc_4558;
wire uc_4559;
wire uc_4560;
wire uc_4561;
wire uc_4562;
wire uc_4563;
wire uc_4564;
wire uc_4565;
wire uc_4566;
wire uc_4567;
wire uc_4568;
wire uc_4569;
wire uc_4570;
wire uc_4571;
wire uc_4572;
wire uc_4573;
wire uc_4574;
wire uc_4575;
wire uc_4576;
wire uc_4577;
wire uc_4578;
wire uc_4579;
wire uc_4580;
wire uc_4581;
wire uc_4582;
wire uc_4583;
wire uc_4584;
wire uc_4585;
wire uc_4586;
wire uc_4587;
wire uc_4588;
wire uc_4589;
wire uc_4590;
wire uc_4591;
wire uc_4592;
wire uc_4593;
wire uc_4594;
wire uc_4595;
wire uc_4596;
wire uc_4597;
wire uc_4598;
wire uc_4599;
wire uc_4600;
wire uc_4601;
wire uc_4602;
wire uc_4603;
wire uc_4604;
wire uc_4605;
wire uc_4606;
wire uc_4607;
wire uc_4608;
wire uc_4609;
wire uc_4610;
wire uc_4611;
wire uc_4612;
wire uc_4613;
wire uc_4614;
wire uc_4615;
wire uc_4616;
wire uc_4617;
wire uc_4618;
wire uc_4619;
wire uc_4620;
wire uc_4621;
wire uc_4622;
wire uc_4623;
wire uc_4624;
wire uc_4625;
wire uc_4626;
wire uc_4627;
wire uc_4628;
wire uc_4629;
wire uc_4630;
wire uc_4631;
wire uc_4632;
wire uc_4633;
wire uc_4634;
wire uc_4635;
wire uc_4636;
wire uc_4637;
wire uc_4638;
wire uc_4639;
wire uc_4640;
wire uc_4641;
wire uc_4642;
wire uc_4643;
wire uc_4644;
wire uc_4645;
wire uc_4646;
wire uc_4647;
wire uc_4648;
wire uc_4649;
wire uc_4650;
wire uc_4651;
wire uc_4652;
wire uc_4653;
wire uc_4654;
wire uc_4655;
wire uc_4656;
wire uc_4657;
wire uc_4658;
wire uc_4659;
wire uc_4660;
wire uc_4661;
wire uc_4662;
wire uc_4663;
wire uc_4664;
wire uc_4665;
wire uc_4666;
wire uc_4667;
wire uc_4668;
wire uc_4669;
wire uc_4670;
wire uc_4671;
wire uc_4672;
wire uc_4673;
wire uc_4674;
wire uc_4675;
wire uc_4676;
wire uc_4677;
wire uc_4678;
wire uc_4679;
wire uc_4680;
wire uc_4681;
wire uc_4682;
wire uc_4683;
wire uc_4684;
wire uc_4685;
wire uc_4686;
wire uc_4687;
wire uc_4688;
wire uc_4689;
wire uc_4690;
wire uc_4691;
wire uc_4692;
wire uc_4693;
wire uc_4694;
wire uc_4695;
wire uc_4696;
wire uc_4697;
wire uc_4698;
wire uc_4699;
wire uc_4700;
wire uc_4701;
wire uc_4702;
wire uc_4703;
wire uc_4704;
wire uc_4705;
wire uc_4706;
wire uc_4707;
wire uc_4708;
wire uc_4709;
wire uc_4710;
wire uc_4711;
wire uc_4712;
wire uc_4713;
wire uc_4714;
wire uc_4715;
wire uc_4716;
wire uc_4717;
wire uc_4718;
wire uc_4719;
wire uc_4720;
wire uc_4721;
wire uc_4722;
wire uc_4723;
wire uc_4724;
wire uc_4725;
wire uc_4726;
wire uc_4727;
wire uc_4728;
wire uc_4729;
wire uc_4730;
wire uc_4731;
wire uc_4732;
wire uc_4733;
wire uc_4734;
wire uc_4735;
wire uc_4736;
wire uc_4737;
wire uc_4738;
wire uc_4739;
wire uc_4740;
wire uc_4741;
wire uc_4742;
wire uc_4743;
wire uc_4744;
wire uc_4745;
wire uc_4746;
wire uc_4747;
wire uc_4748;
wire uc_4749;
wire uc_4750;
wire uc_4751;
wire uc_4752;
wire uc_4753;
wire uc_4754;
wire uc_4755;
wire uc_4756;
wire uc_4757;
wire uc_4758;
wire uc_4759;
wire uc_4760;
wire uc_4761;
wire uc_4762;
wire uc_4763;
wire uc_4764;
wire uc_4765;
wire uc_4766;
wire uc_4767;
wire uc_4768;
wire uc_4769;
wire uc_4770;
wire uc_4771;
wire uc_4772;
wire uc_4773;
wire uc_4774;
wire uc_4775;
wire uc_4776;
wire uc_4777;
wire uc_4778;
wire uc_4779;
wire uc_4780;
wire uc_4781;
wire uc_4782;
wire uc_4783;
wire uc_4784;
wire uc_4785;
wire uc_4786;
wire uc_4787;
wire uc_4788;
wire uc_4789;
wire uc_4790;
wire uc_4791;
wire uc_4792;
wire uc_4793;
wire uc_4794;
wire uc_4795;
wire uc_4796;
wire uc_4797;
wire uc_4798;
wire uc_4799;
wire uc_4800;
wire uc_4801;
wire uc_4802;
wire uc_4803;
wire uc_4804;
wire uc_4805;
wire uc_4806;
wire uc_4807;
wire uc_4808;
wire uc_4809;
wire uc_4810;
wire uc_4811;
wire uc_4812;
wire uc_4813;
wire uc_4814;
wire uc_4815;
wire uc_4816;
wire uc_4817;
wire uc_4818;
wire uc_4819;
wire uc_4820;
wire uc_4821;
wire uc_4822;
wire uc_4823;
wire uc_4824;
wire uc_4825;
wire uc_4826;
wire uc_4827;
wire uc_4828;
wire uc_4829;
wire uc_4830;
wire uc_4831;
wire uc_4832;
wire uc_4833;
wire uc_4834;
wire uc_4835;
wire uc_4836;
wire uc_4837;
wire uc_4838;
wire uc_4839;
wire uc_4840;


RCA64 ripple_adder (.sum ({out[63], out[62], out[61], out[60], out[59], out[58], 
    out[57], out[56], out[55], out[54], out[53], out[52], out[51], out[50], out[49], 
    out[48], out[47], out[46], out[45], out[44], out[43], out[42], out[41], out[40], 
    out[39], out[38], out[37], out[36], out[35], out[34], out[33], out[32], out[31], 
    out[30], out[29], out[28], out[27], out[26], out[25], out[24], out[23], out[22], 
    out[21], out[20], out[19], out[18], out[17], out[16], out[15], out[14], out[13], 
    out[12], out[11], out[10], uc_4831, uc_4832, uc_4833, uc_4834, uc_4835, uc_4836, 
    uc_4837, uc_4838, uc_4839, uc_4840}), .A ({\sums[30][63] , \sums[30][62] , \sums[30][61] , 
    \sums[30][60] , \sums[30][59] , \sums[30][58] , \sums[30][57] , \sums[30][56] , 
    \sums[30][55] , \sums[30][54] , \sums[30][53] , \sums[30][52] , \sums[30][51] , 
    \sums[30][50] , \sums[30][49] , \sums[30][48] , \sums[30][47] , \sums[30][46] , 
    \sums[30][45] , \sums[30][44] , \sums[30][43] , \sums[30][42] , \sums[30][41] , 
    \sums[30][40] , \sums[30][39] , \sums[30][38] , \sums[30][37] , \sums[30][36] , 
    \sums[30][35] , \sums[30][34] , \sums[30][33] , \sums[30][32] , \sums[30][31] , 
    \sums[30][30] , \sums[30][29] , \sums[30][28] , \sums[30][27] , \sums[30][26] , 
    \sums[30][25] , \sums[30][24] , \sums[30][23] , \sums[30][22] , \sums[30][21] , 
    \sums[30][20] , \sums[30][19] , \sums[30][18] , \sums[30][17] , \sums[30][16] , 
    \sums[30][15] , \sums[30][14] , \sums[30][13] , \sums[30][12] , \sums[30][11] , 
    \sums[30][10] , uc_4811, uc_4812, uc_4813, uc_4814, uc_4815, uc_4816, uc_4817, 
    uc_4818, uc_4819, uc_4820}), .B ({\couts[30][63] , \couts[30][62] , \couts[30][61] , 
    \couts[30][60] , \couts[30][59] , \couts[30][58] , \couts[30][57] , \couts[30][56] , 
    \couts[30][55] , \couts[30][54] , \couts[30][53] , \couts[30][52] , \couts[30][51] , 
    \couts[30][50] , \couts[30][49] , \couts[30][48] , \couts[30][47] , \couts[30][46] , 
    \couts[30][45] , \couts[30][44] , \couts[30][43] , \couts[30][42] , \couts[30][41] , 
    \couts[30][40] , \couts[30][39] , \couts[30][38] , \couts[30][37] , \couts[30][36] , 
    \couts[30][35] , \couts[30][34] , \couts[30][33] , \couts[30][32] , \couts[30][31] , 
    \couts[30][30] , \couts[30][29] , \couts[30][28] , \couts[30][27] , \couts[30][26] , 
    \couts[30][25] , \couts[30][24] , \couts[30][23] , \couts[30][22] , \couts[30][21] , 
    \couts[30][20] , \couts[30][19] , \couts[30][18] , \couts[30][17] , \couts[30][16] , 
    \couts[30][15] , \couts[30][14] , \couts[30][13] , \couts[30][12] , \couts[30][11] , 
    \couts[30][10] , uc_4821, uc_4822, uc_4823, uc_4824, uc_4825, uc_4826, uc_4827, 
    uc_4828, uc_4829, uc_4830}));
CSA CSA30 (.u ({\sums[30][63] , \sums[30][62] , \sums[30][61] , \sums[30][60] , \sums[30][59] , 
    \sums[30][58] , \sums[30][57] , \sums[30][56] , \sums[30][55] , \sums[30][54] , 
    \sums[30][53] , \sums[30][52] , \sums[30][51] , \sums[30][50] , \sums[30][49] , 
    \sums[30][48] , \sums[30][47] , \sums[30][46] , \sums[30][45] , \sums[30][44] , 
    \sums[30][43] , \sums[30][42] , \sums[30][41] , \sums[30][40] , \sums[30][39] , 
    \sums[30][38] , \sums[30][37] , \sums[30][36] , \sums[30][35] , \sums[30][34] , 
    \sums[30][33] , \sums[30][32] , \sums[30][31] , \sums[30][30] , \sums[30][29] , 
    \sums[30][28] , \sums[30][27] , \sums[30][26] , \sums[30][25] , \sums[30][24] , 
    \sums[30][23] , \sums[30][22] , \sums[30][21] , \sums[30][20] , \sums[30][19] , 
    \sums[30][18] , \sums[30][17] , \sums[30][16] , \sums[30][15] , \sums[30][14] , 
    \sums[30][13] , \sums[30][12] , \sums[30][11] , \sums[30][10] , out[9], uc_4792, 
    uc_4793, uc_4794, uc_4795, uc_4796, uc_4797, uc_4798, uc_4799, uc_4800}), .v ({
    \couts[30][63] , \couts[30][62] , \couts[30][61] , \couts[30][60] , \couts[30][59] , 
    \couts[30][58] , \couts[30][57] , \couts[30][56] , \couts[30][55] , \couts[30][54] , 
    \couts[30][53] , \couts[30][52] , \couts[30][51] , \couts[30][50] , \couts[30][49] , 
    \couts[30][48] , \couts[30][47] , \couts[30][46] , \couts[30][45] , \couts[30][44] , 
    \couts[30][43] , \couts[30][42] , \couts[30][41] , \couts[30][40] , \couts[30][39] , 
    \couts[30][38] , \couts[30][37] , \couts[30][36] , \couts[30][35] , \couts[30][34] , 
    \couts[30][33] , \couts[30][32] , \couts[30][31] , \couts[30][30] , \couts[30][29] , 
    \couts[30][28] , \couts[30][27] , \couts[30][26] , \couts[30][25] , \couts[30][24] , 
    \couts[30][23] , \couts[30][22] , \couts[30][21] , \couts[30][20] , \couts[30][19] , 
    \couts[30][18] , \couts[30][17] , \couts[30][16] , \couts[30][15] , \couts[30][14] , 
    \couts[30][13] , \couts[30][12] , \couts[30][11] , \couts[30][10] , uc_4801, 
    uc_4802, uc_4803, uc_4804, uc_4805, uc_4806, uc_4807, uc_4808, uc_4809, uc_4810})
    , .x ({\couts[29][63] , \couts[29][62] , \couts[29][61] , \couts[29][60] , \couts[29][59] , 
    \couts[29][58] , \couts[29][57] , \couts[29][56] , \couts[29][55] , \couts[29][54] , 
    \couts[29][53] , \couts[29][52] , \couts[29][51] , \couts[29][50] , \couts[29][49] , 
    \couts[29][48] , \couts[29][47] , \couts[29][46] , \couts[29][45] , \couts[29][44] , 
    \couts[29][43] , \couts[29][42] , \couts[29][41] , \couts[29][40] , \couts[29][39] , 
    \couts[29][38] , \couts[29][37] , \couts[29][36] , \couts[29][35] , \couts[29][34] , 
    \couts[29][33] , \couts[29][32] , \couts[29][31] , \couts[29][30] , \couts[29][29] , 
    \couts[29][28] , \couts[29][27] , \couts[29][26] , \couts[29][25] , \couts[29][24] , 
    \couts[29][23] , \couts[29][22] , \couts[29][21] , \couts[29][20] , \couts[29][19] , 
    \couts[29][18] , \couts[29][17] , \couts[29][16] , \couts[29][15] , \couts[29][14] , 
    \couts[29][13] , \couts[29][12] , \couts[29][11] , \couts[29][10] , \couts[29][9] , 
    uc_4711, uc_4712, uc_4713, uc_4714, uc_4715, uc_4716, uc_4717, uc_4718, uc_4719})
    , .y ({\sums[29][63] , \sums[29][62] , \sums[29][61] , \sums[29][60] , \sums[29][59] , 
    \sums[29][58] , \sums[29][57] , \sums[29][56] , \sums[29][55] , \sums[29][54] , 
    \sums[29][53] , \sums[29][52] , \sums[29][51] , \sums[29][50] , \sums[29][49] , 
    \sums[29][48] , \sums[29][47] , \sums[29][46] , \sums[29][45] , \sums[29][44] , 
    \sums[29][43] , \sums[29][42] , \sums[29][41] , \sums[29][40] , \sums[29][39] , 
    \sums[29][38] , \sums[29][37] , \sums[29][36] , \sums[29][35] , \sums[29][34] , 
    \sums[29][33] , \sums[29][32] , \sums[29][31] , \sums[29][30] , \sums[29][29] , 
    \sums[29][28] , \sums[29][27] , \sums[29][26] , \sums[29][25] , \sums[29][24] , 
    \sums[29][23] , \sums[29][22] , \sums[29][21] , \sums[29][20] , \sums[29][19] , 
    \sums[29][18] , \sums[29][17] , \sums[29][16] , \sums[29][15] , \sums[29][14] , 
    \sums[29][13] , \sums[29][12] , \sums[29][11] , \sums[29][10] , \sums[29][9] , 
    uc_4720, uc_4721, uc_4722, uc_4723, uc_4724, uc_4725, uc_4726, uc_4727, uc_4728})
    , .z ({uc_4729, uc_4730, uc_4731, uc_4732, uc_4733, uc_4734, uc_4735, uc_4736, 
    uc_4737, uc_4738, uc_4739, uc_4740, uc_4741, uc_4742, uc_4743, uc_4744, uc_4745, 
    uc_4746, uc_4747, uc_4748, uc_4749, uc_4750, uc_4751, uc_4752, uc_4753, uc_4754, 
    uc_4755, uc_4756, uc_4757, uc_4758, uc_4759, uc_4760, x[31], uc_4761, uc_4762, 
    uc_4763, uc_4764, uc_4765, uc_4766, uc_4767, uc_4768, uc_4769, uc_4770, uc_4771, 
    uc_4772, uc_4773, uc_4774, uc_4775, uc_4776, uc_4777, uc_4778, uc_4779, uc_4780, 
    uc_4781, uc_4782, uc_4783, uc_4784, uc_4785, uc_4786, uc_4787, uc_4788, uc_4789, 
    uc_4790, uc_4791}));
CSA__5_212 CSA29 (.u ({\sums[29][63] , \sums[29][62] , \sums[29][61] , \sums[29][60] , 
    \sums[29][59] , \sums[29][58] , \sums[29][57] , \sums[29][56] , \sums[29][55] , 
    \sums[29][54] , \sums[29][53] , \sums[29][52] , \sums[29][51] , \sums[29][50] , 
    \sums[29][49] , \sums[29][48] , \sums[29][47] , \sums[29][46] , \sums[29][45] , 
    \sums[29][44] , \sums[29][43] , \sums[29][42] , \sums[29][41] , \sums[29][40] , 
    \sums[29][39] , \sums[29][38] , \sums[29][37] , \sums[29][36] , \sums[29][35] , 
    \sums[29][34] , \sums[29][33] , \sums[29][32] , \sums[29][31] , \sums[29][30] , 
    \sums[29][29] , \sums[29][28] , \sums[29][27] , \sums[29][26] , \sums[29][25] , 
    \sums[29][24] , \sums[29][23] , \sums[29][22] , \sums[29][21] , \sums[29][20] , 
    \sums[29][19] , \sums[29][18] , \sums[29][17] , \sums[29][16] , \sums[29][15] , 
    \sums[29][14] , \sums[29][13] , \sums[29][12] , \sums[29][11] , \sums[29][10] , 
    \sums[29][9] , out[8], uc_4694, uc_4695, uc_4696, uc_4697, uc_4698, uc_4699, 
    uc_4700, uc_4701}), .v ({\couts[29][63] , \couts[29][62] , \couts[29][61] , \couts[29][60] , 
    \couts[29][59] , \couts[29][58] , \couts[29][57] , \couts[29][56] , \couts[29][55] , 
    \couts[29][54] , \couts[29][53] , \couts[29][52] , \couts[29][51] , \couts[29][50] , 
    \couts[29][49] , \couts[29][48] , \couts[29][47] , \couts[29][46] , \couts[29][45] , 
    \couts[29][44] , \couts[29][43] , \couts[29][42] , \couts[29][41] , \couts[29][40] , 
    \couts[29][39] , \couts[29][38] , \couts[29][37] , \couts[29][36] , \couts[29][35] , 
    \couts[29][34] , \couts[29][33] , \couts[29][32] , \couts[29][31] , \couts[29][30] , 
    \couts[29][29] , \couts[29][28] , \couts[29][27] , \couts[29][26] , \couts[29][25] , 
    \couts[29][24] , \couts[29][23] , \couts[29][22] , \couts[29][21] , \couts[29][20] , 
    \couts[29][19] , \couts[29][18] , \couts[29][17] , \couts[29][16] , \couts[29][15] , 
    \couts[29][14] , \couts[29][13] , \couts[29][12] , \couts[29][11] , \couts[29][10] , 
    \couts[29][9] , uc_4702, uc_4703, uc_4704, uc_4705, uc_4706, uc_4707, uc_4708, 
    uc_4709, uc_4710}), .x ({\couts[28][63] , \couts[28][62] , \couts[28][61] , \couts[28][60] , 
    \couts[28][59] , \couts[28][58] , \couts[28][57] , \couts[28][56] , \couts[28][55] , 
    \couts[28][54] , \couts[28][53] , \couts[28][52] , \couts[28][51] , \couts[28][50] , 
    \couts[28][49] , \couts[28][48] , \couts[28][47] , \couts[28][46] , \couts[28][45] , 
    \couts[28][44] , \couts[28][43] , \couts[28][42] , \couts[28][41] , \couts[28][40] , 
    \couts[28][39] , \couts[28][38] , \couts[28][37] , \couts[28][36] , \couts[28][35] , 
    \couts[28][34] , \couts[28][33] , \couts[28][32] , \couts[28][31] , \couts[28][30] , 
    \couts[28][29] , \couts[28][28] , \couts[28][27] , \couts[28][26] , \couts[28][25] , 
    \couts[28][24] , \couts[28][23] , \couts[28][22] , \couts[28][21] , \couts[28][20] , 
    \couts[28][19] , \couts[28][18] , \couts[28][17] , \couts[28][16] , \couts[28][15] , 
    \couts[28][14] , \couts[28][13] , \couts[28][12] , \couts[28][11] , \couts[28][10] , 
    \couts[28][9] , \couts[28][8] , uc_4647, uc_4648, uc_4649, uc_4650, uc_4651, 
    uc_4652, uc_4653, uc_4654}), .y ({\sums[28][63] , \sums[28][62] , \sums[28][61] , 
    \sums[28][60] , \sums[28][59] , \sums[28][58] , \sums[28][57] , \sums[28][56] , 
    \sums[28][55] , \sums[28][54] , \sums[28][53] , \sums[28][52] , \sums[28][51] , 
    \sums[28][50] , \sums[28][49] , \sums[28][48] , \sums[28][47] , \sums[28][46] , 
    \sums[28][45] , \sums[28][44] , \sums[28][43] , \sums[28][42] , \sums[28][41] , 
    \sums[28][40] , \sums[28][39] , \sums[28][38] , \sums[28][37] , \sums[28][36] , 
    \sums[28][35] , \sums[28][34] , \sums[28][33] , \sums[28][32] , \sums[28][31] , 
    \sums[28][30] , \sums[28][29] , \sums[28][28] , \sums[28][27] , \sums[28][26] , 
    \sums[28][25] , \sums[28][24] , \sums[28][23] , \sums[28][22] , \sums[28][21] , 
    \sums[28][20] , \sums[28][19] , \sums[28][18] , \sums[28][17] , \sums[28][16] , 
    \sums[28][15] , \sums[28][14] , \sums[28][13] , \sums[28][12] , \sums[28][11] , 
    \sums[28][10] , \sums[28][9] , \sums[28][8] , uc_4655, uc_4656, uc_4657, uc_4658, 
    uc_4659, uc_4660, uc_4661, uc_4662}), .z ({\couts[21][63] , \couts[21][62] , 
    \couts[21][61] , \couts[21][60] , \couts[21][59] , \couts[21][58] , \couts[21][57] , 
    \couts[21][56] , \couts[21][55] , \couts[21][54] , \couts[21][53] , \couts[21][52] , 
    \couts[21][51] , \couts[21][50] , \couts[21][49] , \couts[21][48] , \couts[21][47] , 
    \couts[21][46] , \couts[21][45] , \couts[21][44] , \couts[21][43] , \couts[21][42] , 
    \couts[21][41] , \couts[21][40] , \couts[21][39] , \couts[21][38] , \couts[21][37] , 
    \couts[21][36] , \couts[21][35] , \couts[21][34] , \couts[21][33] , \couts[21][32] , 
    \couts[21][31] , uc_4663, uc_4664, uc_4665, uc_4666, uc_4667, uc_4668, uc_4669, 
    uc_4670, uc_4671, uc_4672, uc_4673, uc_4674, uc_4675, uc_4676, uc_4677, uc_4678, 
    uc_4679, uc_4680, uc_4681, uc_4682, uc_4683, uc_4684, uc_4685, uc_4686, uc_4687, 
    uc_4688, uc_4689, uc_4690, uc_4691, uc_4692, uc_4693}));
CSA__5_209 CSA28 (.u ({\sums[28][63] , \sums[28][62] , \sums[28][61] , \sums[28][60] , 
    \sums[28][59] , \sums[28][58] , \sums[28][57] , \sums[28][56] , \sums[28][55] , 
    \sums[28][54] , \sums[28][53] , \sums[28][52] , \sums[28][51] , \sums[28][50] , 
    \sums[28][49] , \sums[28][48] , \sums[28][47] , \sums[28][46] , \sums[28][45] , 
    \sums[28][44] , \sums[28][43] , \sums[28][42] , \sums[28][41] , \sums[28][40] , 
    \sums[28][39] , \sums[28][38] , \sums[28][37] , \sums[28][36] , \sums[28][35] , 
    \sums[28][34] , \sums[28][33] , \sums[28][32] , \sums[28][31] , \sums[28][30] , 
    \sums[28][29] , \sums[28][28] , \sums[28][27] , \sums[28][26] , \sums[28][25] , 
    \sums[28][24] , \sums[28][23] , \sums[28][22] , \sums[28][21] , \sums[28][20] , 
    \sums[28][19] , \sums[28][18] , \sums[28][17] , \sums[28][16] , \sums[28][15] , 
    \sums[28][14] , \sums[28][13] , \sums[28][12] , \sums[28][11] , \sums[28][10] , 
    \sums[28][9] , \sums[28][8] , out[7], uc_4632, uc_4633, uc_4634, uc_4635, uc_4636, 
    uc_4637, uc_4638}), .v ({\couts[28][63] , \couts[28][62] , \couts[28][61] , \couts[28][60] , 
    \couts[28][59] , \couts[28][58] , \couts[28][57] , \couts[28][56] , \couts[28][55] , 
    \couts[28][54] , \couts[28][53] , \couts[28][52] , \couts[28][51] , \couts[28][50] , 
    \couts[28][49] , \couts[28][48] , \couts[28][47] , \couts[28][46] , \couts[28][45] , 
    \couts[28][44] , \couts[28][43] , \couts[28][42] , \couts[28][41] , \couts[28][40] , 
    \couts[28][39] , \couts[28][38] , \couts[28][37] , \couts[28][36] , \couts[28][35] , 
    \couts[28][34] , \couts[28][33] , \couts[28][32] , \couts[28][31] , \couts[28][30] , 
    \couts[28][29] , \couts[28][28] , \couts[28][27] , \couts[28][26] , \couts[28][25] , 
    \couts[28][24] , \couts[28][23] , \couts[28][22] , \couts[28][21] , \couts[28][20] , 
    \couts[28][19] , \couts[28][18] , \couts[28][17] , \couts[28][16] , \couts[28][15] , 
    \couts[28][14] , \couts[28][13] , \couts[28][12] , \couts[28][11] , \couts[28][10] , 
    \couts[28][9] , \couts[28][8] , uc_4639, uc_4640, uc_4641, uc_4642, uc_4643, 
    uc_4644, uc_4645, uc_4646}), .x ({\couts[27][63] , \couts[27][62] , \couts[27][61] , 
    \couts[27][60] , \couts[27][59] , \couts[27][58] , \couts[27][57] , \couts[27][56] , 
    \couts[27][55] , \couts[27][54] , \couts[27][53] , \couts[27][52] , \couts[27][51] , 
    \couts[27][50] , \couts[27][49] , \couts[27][48] , \couts[27][47] , \couts[27][46] , 
    \couts[27][45] , \couts[27][44] , \couts[27][43] , \couts[27][42] , \couts[27][41] , 
    \couts[27][40] , \couts[27][39] , \couts[27][38] , \couts[27][37] , \couts[27][36] , 
    \couts[27][35] , \couts[27][34] , \couts[27][33] , \couts[27][32] , \couts[27][31] , 
    \couts[27][30] , \couts[27][29] , \couts[27][28] , \couts[27][27] , \couts[27][26] , 
    \couts[27][25] , \couts[27][24] , \couts[27][23] , \couts[27][22] , \couts[27][21] , 
    \couts[27][20] , \couts[27][19] , \couts[27][18] , \couts[27][17] , \couts[27][16] , 
    \couts[27][15] , \couts[27][14] , \couts[27][13] , \couts[27][12] , \couts[27][11] , 
    \couts[27][10] , \couts[27][9] , \couts[27][8] , \couts[27][7] , uc_4596, uc_4597, 
    uc_4598, uc_4599, uc_4600, uc_4601, uc_4602}), .y ({\sums[27][63] , \sums[27][62] , 
    \sums[27][61] , \sums[27][60] , \sums[27][59] , \sums[27][58] , \sums[27][57] , 
    \sums[27][56] , \sums[27][55] , \sums[27][54] , \sums[27][53] , \sums[27][52] , 
    \sums[27][51] , \sums[27][50] , \sums[27][49] , \sums[27][48] , \sums[27][47] , 
    \sums[27][46] , \sums[27][45] , \sums[27][44] , \sums[27][43] , \sums[27][42] , 
    \sums[27][41] , \sums[27][40] , \sums[27][39] , \sums[27][38] , \sums[27][37] , 
    \sums[27][36] , \sums[27][35] , \sums[27][34] , \sums[27][33] , \sums[27][32] , 
    \sums[27][31] , \sums[27][30] , \sums[27][29] , \sums[27][28] , \sums[27][27] , 
    \sums[27][26] , \sums[27][25] , \sums[27][24] , \sums[27][23] , \sums[27][22] , 
    \sums[27][21] , \sums[27][20] , \sums[27][19] , \sums[27][18] , \sums[27][17] , 
    \sums[27][16] , \sums[27][15] , \sums[27][14] , \sums[27][13] , \sums[27][12] , 
    \sums[27][11] , \sums[27][10] , \sums[27][9] , \sums[27][8] , \sums[27][7] , 
    uc_4603, uc_4604, uc_4605, uc_4606, uc_4607, uc_4608, uc_4609}), .z ({\couts[26][63] , 
    \couts[26][62] , \couts[26][61] , \couts[26][60] , \couts[26][59] , \couts[26][58] , 
    \couts[26][57] , \couts[26][56] , \couts[26][55] , \couts[26][54] , \couts[26][53] , 
    \couts[26][52] , \couts[26][51] , \couts[26][50] , \couts[26][49] , \couts[26][48] , 
    \couts[26][47] , \couts[26][46] , \couts[26][45] , \couts[26][44] , \couts[26][43] , 
    \couts[26][42] , \couts[26][41] , \couts[26][40] , \couts[26][39] , \couts[26][38] , 
    \couts[26][37] , \couts[26][36] , \couts[26][35] , \couts[26][34] , \couts[26][33] , 
    \couts[26][32] , \couts[26][31] , \couts[26][30] , \couts[26][29] , \couts[26][28] , 
    \couts[26][27] , \couts[26][26] , \couts[26][25] , \couts[26][24] , \couts[26][23] , 
    \couts[26][22] , uc_4610, uc_4611, uc_4612, uc_4613, uc_4614, uc_4615, uc_4616, 
    uc_4617, uc_4618, uc_4619, uc_4620, uc_4621, uc_4622, uc_4623, uc_4624, uc_4625, 
    uc_4626, uc_4627, uc_4628, uc_4629, uc_4630, uc_4631}));
CSA__5_206 CSA27 (.u ({\sums[27][63] , \sums[27][62] , \sums[27][61] , \sums[27][60] , 
    \sums[27][59] , \sums[27][58] , \sums[27][57] , \sums[27][56] , \sums[27][55] , 
    \sums[27][54] , \sums[27][53] , \sums[27][52] , \sums[27][51] , \sums[27][50] , 
    \sums[27][49] , \sums[27][48] , \sums[27][47] , \sums[27][46] , \sums[27][45] , 
    \sums[27][44] , \sums[27][43] , \sums[27][42] , \sums[27][41] , \sums[27][40] , 
    \sums[27][39] , \sums[27][38] , \sums[27][37] , \sums[27][36] , \sums[27][35] , 
    \sums[27][34] , \sums[27][33] , \sums[27][32] , \sums[27][31] , \sums[27][30] , 
    \sums[27][29] , \sums[27][28] , \sums[27][27] , \sums[27][26] , \sums[27][25] , 
    \sums[27][24] , \sums[27][23] , \sums[27][22] , \sums[27][21] , \sums[27][20] , 
    \sums[27][19] , \sums[27][18] , \sums[27][17] , \sums[27][16] , \sums[27][15] , 
    \sums[27][14] , \sums[27][13] , \sums[27][12] , \sums[27][11] , \sums[27][10] , 
    \sums[27][9] , \sums[27][8] , \sums[27][7] , out[6], uc_4583, uc_4584, uc_4585, 
    uc_4586, uc_4587, uc_4588}), .v ({\couts[27][63] , \couts[27][62] , \couts[27][61] , 
    \couts[27][60] , \couts[27][59] , \couts[27][58] , \couts[27][57] , \couts[27][56] , 
    \couts[27][55] , \couts[27][54] , \couts[27][53] , \couts[27][52] , \couts[27][51] , 
    \couts[27][50] , \couts[27][49] , \couts[27][48] , \couts[27][47] , \couts[27][46] , 
    \couts[27][45] , \couts[27][44] , \couts[27][43] , \couts[27][42] , \couts[27][41] , 
    \couts[27][40] , \couts[27][39] , \couts[27][38] , \couts[27][37] , \couts[27][36] , 
    \couts[27][35] , \couts[27][34] , \couts[27][33] , \couts[27][32] , \couts[27][31] , 
    \couts[27][30] , \couts[27][29] , \couts[27][28] , \couts[27][27] , \couts[27][26] , 
    \couts[27][25] , \couts[27][24] , \couts[27][23] , \couts[27][22] , \couts[27][21] , 
    \couts[27][20] , \couts[27][19] , \couts[27][18] , \couts[27][17] , \couts[27][16] , 
    \couts[27][15] , \couts[27][14] , \couts[27][13] , \couts[27][12] , \couts[27][11] , 
    \couts[27][10] , \couts[27][9] , \couts[27][8] , \couts[27][7] , uc_4589, uc_4590, 
    uc_4591, uc_4592, uc_4593, uc_4594, uc_4595}), .x ({\sums[25][63] , \sums[25][62] , 
    \sums[25][61] , \sums[25][60] , \sums[25][59] , \sums[25][58] , \sums[25][57] , 
    \sums[25][56] , \sums[25][55] , \sums[25][54] , \sums[25][53] , \sums[25][52] , 
    \sums[25][51] , \sums[25][50] , \sums[25][49] , \sums[25][48] , \sums[25][47] , 
    \sums[25][46] , \sums[25][45] , \sums[25][44] , \sums[25][43] , \sums[25][42] , 
    \sums[25][41] , \sums[25][40] , \sums[25][39] , \sums[25][38] , \sums[25][37] , 
    \sums[25][36] , \sums[25][35] , \sums[25][34] , \sums[25][33] , \sums[25][32] , 
    \sums[25][31] , \sums[25][30] , \sums[25][29] , \sums[25][28] , \sums[25][27] , 
    \sums[25][26] , \sums[25][25] , \sums[25][24] , \sums[25][23] , \sums[25][22] , 
    \sums[25][21] , \sums[25][20] , \sums[25][19] , \sums[25][18] , \sums[25][17] , 
    \sums[25][16] , \sums[25][15] , \sums[25][14] , \sums[25][13] , \sums[25][12] , 
    \sums[25][11] , \sums[25][10] , \sums[25][9] , \sums[25][8] , \sums[25][7] , 
    \sums[25][6] , uc_4556, uc_4557, uc_4558, uc_4559, uc_4560, uc_4561}), .y ({\couts[25][63] , 
    \couts[25][62] , \couts[25][61] , \couts[25][60] , \couts[25][59] , \couts[25][58] , 
    \couts[25][57] , \couts[25][56] , \couts[25][55] , \couts[25][54] , \couts[25][53] , 
    \couts[25][52] , \couts[25][51] , \couts[25][50] , \couts[25][49] , \couts[25][48] , 
    \couts[25][47] , \couts[25][46] , \couts[25][45] , \couts[25][44] , \couts[25][43] , 
    \couts[25][42] , \couts[25][41] , \couts[25][40] , \couts[25][39] , \couts[25][38] , 
    \couts[25][37] , \couts[25][36] , \couts[25][35] , \couts[25][34] , \couts[25][33] , 
    \couts[25][32] , \couts[25][31] , \couts[25][30] , \couts[25][29] , \couts[25][28] , 
    \couts[25][27] , \couts[25][26] , \couts[25][25] , \couts[25][24] , \couts[25][23] , 
    \couts[25][22] , \couts[25][21] , \couts[25][20] , \couts[25][19] , \couts[25][18] , 
    \couts[25][17] , \couts[25][16] , \couts[25][15] , \couts[25][14] , \couts[25][13] , 
    \couts[25][12] , \couts[25][11] , \couts[25][10] , \couts[25][9] , \couts[25][8] , 
    \couts[25][7] , \couts[25][6] , uc_4562, uc_4563, uc_4564, uc_4565, uc_4566, 
    uc_4567}), .z ({\sums[26][63] , \sums[26][62] , \sums[26][61] , \sums[26][60] , 
    \sums[26][59] , \sums[26][58] , \sums[26][57] , \sums[26][56] , \sums[26][55] , 
    \sums[26][54] , \sums[26][53] , \sums[26][52] , \sums[26][51] , \sums[26][50] , 
    \sums[26][49] , \sums[26][48] , \sums[26][47] , \sums[26][46] , \sums[26][45] , 
    \sums[26][44] , \sums[26][43] , \sums[26][42] , \sums[26][41] , \sums[26][40] , 
    \sums[26][39] , \sums[26][38] , \sums[26][37] , \sums[26][36] , \sums[26][35] , 
    \sums[26][34] , \sums[26][33] , \sums[26][32] , \sums[26][31] , \sums[26][30] , 
    \sums[26][29] , \sums[26][28] , \sums[26][27] , \sums[26][26] , \sums[26][25] , 
    \sums[26][24] , \sums[26][23] , \sums[26][22] , \sums[26][21] , \couts[23][20] , 
    \couts[23][19] , \couts[23][18] , \couts[23][17] , \couts[23][16] , \couts[23][15] , 
    uc_4568, uc_4569, uc_4570, uc_4571, uc_4572, uc_4573, uc_4574, uc_4575, uc_4576, 
    uc_4577, uc_4578, uc_4579, uc_4580, uc_4581, uc_4582}));
CSA__5_203 CSA26 (.u ({\sums[26][63] , \sums[26][62] , \sums[26][61] , \sums[26][60] , 
    \sums[26][59] , \sums[26][58] , \sums[26][57] , \sums[26][56] , \sums[26][55] , 
    \sums[26][54] , \sums[26][53] , \sums[26][52] , \sums[26][51] , \sums[26][50] , 
    \sums[26][49] , \sums[26][48] , \sums[26][47] , \sums[26][46] , \sums[26][45] , 
    \sums[26][44] , \sums[26][43] , \sums[26][42] , \sums[26][41] , \sums[26][40] , 
    \sums[26][39] , \sums[26][38] , \sums[26][37] , \sums[26][36] , \sums[26][35] , 
    \sums[26][34] , \sums[26][33] , \sums[26][32] , \sums[26][31] , \sums[26][30] , 
    \sums[26][29] , \sums[26][28] , \sums[26][27] , \sums[26][26] , \sums[26][25] , 
    \sums[26][24] , \sums[26][23] , \sums[26][22] , \sums[26][21] , uc_4513, uc_4514, 
    uc_4515, uc_4516, uc_4517, uc_4518, uc_4519, uc_4520, uc_4521, uc_4522, uc_4523, 
    uc_4524, uc_4525, uc_4526, uc_4527, uc_4528, uc_4529, uc_4530, uc_4531, uc_4532, 
    uc_4533}), .v ({\couts[26][63] , \couts[26][62] , \couts[26][61] , \couts[26][60] , 
    \couts[26][59] , \couts[26][58] , \couts[26][57] , \couts[26][56] , \couts[26][55] , 
    \couts[26][54] , \couts[26][53] , \couts[26][52] , \couts[26][51] , \couts[26][50] , 
    \couts[26][49] , \couts[26][48] , \couts[26][47] , \couts[26][46] , \couts[26][45] , 
    \couts[26][44] , \couts[26][43] , \couts[26][42] , \couts[26][41] , \couts[26][40] , 
    \couts[26][39] , \couts[26][38] , \couts[26][37] , \couts[26][36] , \couts[26][35] , 
    \couts[26][34] , \couts[26][33] , \couts[26][32] , \couts[26][31] , \couts[26][30] , 
    \couts[26][29] , \couts[26][28] , \couts[26][27] , \couts[26][26] , \couts[26][25] , 
    \couts[26][24] , \couts[26][23] , \couts[26][22] , uc_4534, uc_4535, uc_4536, 
    uc_4537, uc_4538, uc_4539, uc_4540, uc_4541, uc_4542, uc_4543, uc_4544, uc_4545, 
    uc_4546, uc_4547, uc_4548, uc_4549, uc_4550, uc_4551, uc_4552, uc_4553, uc_4554, 
    uc_4555}), .x ({\couts[23][63] , \couts[23][62] , \couts[23][61] , \couts[23][60] , 
    \couts[23][59] , \couts[23][58] , \couts[23][57] , \couts[23][56] , \couts[23][55] , 
    \couts[23][54] , \couts[23][53] , \couts[23][52] , \couts[23][51] , \couts[23][50] , 
    \couts[23][49] , \couts[23][48] , \couts[23][47] , \couts[23][46] , \couts[23][45] , 
    \couts[23][44] , \couts[23][43] , \couts[23][42] , \couts[23][41] , \couts[23][40] , 
    \couts[23][39] , \couts[23][38] , \couts[23][37] , \couts[23][36] , \couts[23][35] , 
    \couts[23][34] , \couts[23][33] , \couts[23][32] , \couts[23][31] , \couts[23][30] , 
    \couts[23][29] , \couts[23][28] , \couts[23][27] , \couts[23][26] , \couts[23][25] , 
    \couts[23][24] , \couts[23][23] , \couts[23][22] , \couts[23][21] , uc_4446, 
    uc_4447, uc_4448, uc_4449, uc_4450, uc_4451, uc_4452, uc_4453, uc_4454, uc_4455, 
    uc_4456, uc_4457, uc_4458, uc_4459, uc_4460, uc_4461, uc_4462, uc_4463, uc_4464, 
    uc_4465, uc_4466}), .y ({\sums[24][63] , \sums[24][62] , \sums[24][61] , \sums[24][60] , 
    \sums[24][59] , \sums[24][58] , \sums[24][57] , \sums[24][56] , \sums[24][55] , 
    \sums[24][54] , \sums[24][53] , \sums[24][52] , \sums[24][51] , \sums[24][50] , 
    \sums[24][49] , \sums[24][48] , \sums[24][47] , \sums[24][46] , \sums[24][45] , 
    \sums[24][44] , \sums[24][43] , \sums[24][42] , \sums[24][41] , \sums[24][40] , 
    \sums[24][39] , \sums[24][38] , \sums[24][37] , \sums[24][36] , \sums[24][35] , 
    \sums[24][34] , \sums[24][33] , \sums[24][32] , \sums[24][31] , \sums[24][30] , 
    \sums[24][29] , \sums[24][28] , \sums[24][27] , \sums[24][26] , \sums[24][25] , 
    \sums[24][24] , \sums[20][23] , \sums[20][22] , \sums[20][21] , uc_4467, uc_4468, 
    uc_4469, uc_4470, uc_4471, uc_4472, uc_4473, uc_4474, uc_4475, uc_4476, uc_4477, 
    uc_4478, uc_4479, uc_4480, uc_4481, uc_4482, uc_4483, uc_4484, uc_4485, uc_4486, 
    uc_4487}), .z ({\couts[24][63] , \couts[24][62] , \couts[24][61] , \couts[24][60] , 
    \couts[24][59] , \couts[24][58] , \couts[24][57] , \couts[24][56] , \couts[24][55] , 
    \couts[24][54] , \couts[24][53] , \couts[24][52] , \couts[24][51] , \couts[24][50] , 
    \couts[24][49] , \couts[24][48] , \couts[24][47] , \couts[24][46] , \couts[24][45] , 
    \couts[24][44] , \couts[24][43] , \couts[24][42] , \couts[24][41] , \couts[24][40] , 
    \couts[24][39] , \couts[24][38] , \couts[24][37] , \couts[24][36] , \couts[24][35] , 
    \couts[24][34] , \couts[24][33] , \couts[24][32] , \couts[24][31] , \couts[24][30] , 
    \couts[24][29] , \couts[24][28] , \couts[24][27] , \couts[24][26] , \couts[24][25] , 
    uc_4488, uc_4489, uc_4490, uc_4491, uc_4492, uc_4493, uc_4494, uc_4495, uc_4496, 
    uc_4497, uc_4498, uc_4499, uc_4500, uc_4501, uc_4502, uc_4503, uc_4504, uc_4505, 
    uc_4506, uc_4507, uc_4508, uc_4509, uc_4510, uc_4511, uc_4512}));
CSA__5_200 CSA24 (.u ({\sums[24][63] , \sums[24][62] , \sums[24][61] , \sums[24][60] , 
    \sums[24][59] , \sums[24][58] , \sums[24][57] , \sums[24][56] , \sums[24][55] , 
    \sums[24][54] , \sums[24][53] , \sums[24][52] , \sums[24][51] , \sums[24][50] , 
    \sums[24][49] , \sums[24][48] , \sums[24][47] , \sums[24][46] , \sums[24][45] , 
    \sums[24][44] , \sums[24][43] , \sums[24][42] , \sums[24][41] , \sums[24][40] , 
    \sums[24][39] , \sums[24][38] , \sums[24][37] , \sums[24][36] , \sums[24][35] , 
    \sums[24][34] , \sums[24][33] , \sums[24][32] , \sums[24][31] , \sums[24][30] , 
    \sums[24][29] , \sums[24][28] , \sums[24][27] , \sums[24][26] , \sums[24][25] , 
    \sums[24][24] , uc_4397, uc_4398, uc_4399, uc_4400, uc_4401, uc_4402, uc_4403, 
    uc_4404, uc_4405, uc_4406, uc_4407, uc_4408, uc_4409, uc_4410, uc_4411, uc_4412, 
    uc_4413, uc_4414, uc_4415, uc_4416, uc_4417, uc_4418, uc_4419, uc_4420}), .v ({
    \couts[24][63] , \couts[24][62] , \couts[24][61] , \couts[24][60] , \couts[24][59] , 
    \couts[24][58] , \couts[24][57] , \couts[24][56] , \couts[24][55] , \couts[24][54] , 
    \couts[24][53] , \couts[24][52] , \couts[24][51] , \couts[24][50] , \couts[24][49] , 
    \couts[24][48] , \couts[24][47] , \couts[24][46] , \couts[24][45] , \couts[24][44] , 
    \couts[24][43] , \couts[24][42] , \couts[24][41] , \couts[24][40] , \couts[24][39] , 
    \couts[24][38] , \couts[24][37] , \couts[24][36] , \couts[24][35] , \couts[24][34] , 
    \couts[24][33] , \couts[24][32] , \couts[24][31] , \couts[24][30] , \couts[24][29] , 
    \couts[24][28] , \couts[24][27] , \couts[24][26] , \couts[24][25] , uc_4421, 
    uc_4422, uc_4423, uc_4424, uc_4425, uc_4426, uc_4427, uc_4428, uc_4429, uc_4430, 
    uc_4431, uc_4432, uc_4433, uc_4434, uc_4435, uc_4436, uc_4437, uc_4438, uc_4439, 
    uc_4440, uc_4441, uc_4442, uc_4443, uc_4444, uc_4445}), .x ({\sums[20][59] , 
    \sums[20][59] , \sums[20][59] , \sums[20][59] , \sums[20][59] , \sums[20][58] , 
    \sums[20][57] , \sums[20][56] , \sums[20][55] , \sums[20][54] , \sums[20][53] , 
    \sums[20][52] , \sums[20][51] , \sums[20][50] , \sums[20][49] , \sums[20][48] , 
    \sums[20][47] , \sums[20][46] , \sums[20][45] , \sums[20][44] , \sums[20][43] , 
    \sums[20][42] , \sums[20][41] , \sums[20][40] , \sums[20][39] , \sums[20][38] , 
    \sums[20][37] , \sums[20][36] , \sums[20][35] , \sums[20][34] , \sums[20][33] , 
    \sums[20][32] , \sums[20][31] , \sums[20][30] , \sums[20][29] , \sums[20][28] , 
    \sums[20][27] , \sums[20][26] , \sums[20][25] , \sums[20][24] , uc_4319, uc_4320, 
    uc_4321, uc_4322, uc_4323, uc_4324, uc_4325, uc_4326, uc_4327, uc_4328, uc_4329, 
    uc_4330, uc_4331, uc_4332, uc_4333, uc_4334, uc_4335, uc_4336, uc_4337, uc_4338, 
    uc_4339, uc_4340, uc_4341, uc_4342}), .y ({\couts[20][63] , uc_4343, uc_4344, 
    uc_4345, \couts[20][59] , \couts[20][58] , \couts[20][57] , \couts[20][56] , 
    \couts[20][55] , \couts[20][54] , \couts[20][53] , \couts[20][52] , \couts[20][51] , 
    \couts[20][50] , \couts[20][49] , \couts[20][48] , \couts[20][47] , \couts[20][46] , 
    \couts[20][45] , \couts[20][44] , \couts[20][43] , \couts[20][42] , \couts[20][41] , 
    \couts[20][40] , \couts[20][39] , \couts[20][38] , \couts[20][37] , \couts[20][36] , 
    \couts[20][35] , \couts[20][34] , \couts[20][33] , \couts[20][32] , \couts[20][31] , 
    \couts[20][30] , \couts[20][29] , \couts[20][28] , \couts[20][27] , \couts[20][26] , 
    \couts[20][25] , \couts[20][24] , uc_4346, uc_4347, uc_4348, uc_4349, uc_4350, 
    uc_4351, uc_4352, uc_4353, uc_4354, uc_4355, uc_4356, uc_4357, uc_4358, uc_4359, 
    uc_4360, uc_4361, uc_4362, uc_4363, uc_4364, uc_4365, uc_4366, uc_4367, uc_4368, 
    uc_4369}), .z ({\sums[21][63] , \sums[21][62] , \sums[21][61] , \sums[21][60] , 
    \sums[21][59] , \sums[21][58] , \sums[21][57] , \sums[21][56] , \sums[21][55] , 
    \sums[21][54] , \sums[21][53] , \sums[21][52] , \sums[21][51] , \sums[21][50] , 
    \sums[21][49] , \sums[21][48] , \sums[21][47] , \sums[21][46] , \sums[21][45] , 
    \sums[21][44] , \sums[21][43] , \sums[21][42] , \sums[21][41] , \sums[21][40] , 
    \sums[21][39] , \sums[21][38] , \sums[21][37] , \sums[21][36] , \sums[21][35] , 
    \sums[21][34] , \sums[21][33] , \sums[21][32] , \sums[21][31] , \sums[21][30] , 
    \sums[16][29] , \sums[9][28] , \pp[27][27] , uc_4370, uc_4371, uc_4372, uc_4373, 
    uc_4374, uc_4375, uc_4376, uc_4377, uc_4378, uc_4379, uc_4380, uc_4381, uc_4382, 
    uc_4383, uc_4384, uc_4385, uc_4386, uc_4387, uc_4388, uc_4389, uc_4390, uc_4391, 
    uc_4392, uc_4393, uc_4394, uc_4395, uc_4396}));
CSA__5_197 CSA21 (.u ({\sums[21][63] , \sums[21][62] , \sums[21][61] , \sums[21][60] , 
    \sums[21][59] , \sums[21][58] , \sums[21][57] , \sums[21][56] , \sums[21][55] , 
    \sums[21][54] , \sums[21][53] , \sums[21][52] , \sums[21][51] , \sums[21][50] , 
    \sums[21][49] , \sums[21][48] , \sums[21][47] , \sums[21][46] , \sums[21][45] , 
    \sums[21][44] , \sums[21][43] , \sums[21][42] , \sums[21][41] , \sums[21][40] , 
    \sums[21][39] , \sums[21][38] , \sums[21][37] , \sums[21][36] , \sums[21][35] , 
    \sums[21][34] , \sums[21][33] , \sums[21][32] , \sums[21][31] , \sums[21][30] , 
    uc_4258, uc_4259, uc_4260, uc_4261, uc_4262, uc_4263, uc_4264, uc_4265, uc_4266, 
    uc_4267, uc_4268, uc_4269, uc_4270, uc_4271, uc_4272, uc_4273, uc_4274, uc_4275, 
    uc_4276, uc_4277, uc_4278, uc_4279, uc_4280, uc_4281, uc_4282, uc_4283, uc_4284, 
    uc_4285, uc_4286, uc_4287}), .v ({\couts[21][63] , \couts[21][62] , \couts[21][61] , 
    \couts[21][60] , \couts[21][59] , \couts[21][58] , \couts[21][57] , \couts[21][56] , 
    \couts[21][55] , \couts[21][54] , \couts[21][53] , \couts[21][52] , \couts[21][51] , 
    \couts[21][50] , \couts[21][49] , \couts[21][48] , \couts[21][47] , \couts[21][46] , 
    \couts[21][45] , \couts[21][44] , \couts[21][43] , \couts[21][42] , \couts[21][41] , 
    \couts[21][40] , \couts[21][39] , \couts[21][38] , \couts[21][37] , \couts[21][36] , 
    \couts[21][35] , \couts[21][34] , \couts[21][33] , \couts[21][32] , \couts[21][31] , 
    uc_4288, uc_4289, uc_4290, uc_4291, uc_4292, uc_4293, uc_4294, uc_4295, uc_4296, 
    uc_4297, uc_4298, uc_4299, uc_4300, uc_4301, uc_4302, uc_4303, uc_4304, uc_4305, 
    uc_4306, uc_4307, uc_4308, uc_4309, uc_4310, uc_4311, uc_4312, uc_4313, uc_4314, 
    uc_4315, uc_4316, uc_4317, uc_4318}), .x ({\sums[16][63] , \sums[16][62] , \sums[16][61] , 
    \sums[16][60] , \sums[16][59] , \sums[16][58] , \sums[16][57] , \sums[16][56] , 
    \sums[16][55] , \sums[16][54] , \sums[16][53] , \sums[16][52] , \sums[16][51] , 
    \sums[16][50] , \sums[16][49] , \sums[16][48] , \sums[16][47] , \sums[16][46] , 
    \sums[16][45] , \sums[16][44] , \sums[16][43] , \sums[16][42] , \sums[16][41] , 
    \sums[16][40] , \sums[16][39] , \sums[16][38] , \sums[16][37] , \sums[16][36] , 
    \sums[16][35] , \sums[16][34] , \sums[16][33] , \sums[16][32] , \sums[16][31] , 
    \sums[16][30] , uc_4166, uc_4167, uc_4168, uc_4169, uc_4170, uc_4171, uc_4172, 
    uc_4173, uc_4174, uc_4175, uc_4176, uc_4177, uc_4178, uc_4179, uc_4180, uc_4181, 
    uc_4182, uc_4183, uc_4184, uc_4185, uc_4186, uc_4187, uc_4188, uc_4189, uc_4190, 
    uc_4191, uc_4192, uc_4193, uc_4194, uc_4195}), .y ({\couts[16][63] , \couts[16][62] , 
    \couts[16][61] , \couts[16][60] , \couts[16][59] , \couts[16][58] , \couts[16][57] , 
    \couts[16][56] , \couts[16][55] , \couts[16][54] , \couts[16][53] , \couts[16][52] , 
    \couts[16][51] , \couts[16][50] , \couts[16][49] , \couts[16][48] , \couts[16][47] , 
    \couts[16][46] , \couts[16][45] , \couts[16][44] , \couts[16][43] , \couts[16][42] , 
    \couts[16][41] , \couts[16][40] , \couts[16][39] , \couts[16][38] , \couts[16][37] , 
    \couts[16][36] , \couts[16][35] , \couts[16][34] , \couts[16][33] , \couts[16][32] , 
    \couts[16][31] , \couts[16][30] , uc_4196, uc_4197, uc_4198, uc_4199, uc_4200, 
    uc_4201, uc_4202, uc_4203, uc_4204, uc_4205, uc_4206, uc_4207, uc_4208, uc_4209, 
    uc_4210, uc_4211, uc_4212, uc_4213, uc_4214, uc_4215, uc_4216, uc_4217, uc_4218, 
    uc_4219, uc_4220, uc_4221, uc_4222, uc_4223, uc_4224, uc_4225}), .z ({\pp[31][63] , 
    uc_4226, \pp[31][61] , \pp[31][60] , \pp[31][59] , \pp[31][58] , \pp[31][57] , 
    \pp[31][56] , \pp[31][55] , \pp[31][54] , \pp[31][53] , \pp[31][52] , \pp[31][51] , 
    \pp[31][50] , \pp[31][49] , \pp[31][48] , \pp[31][47] , \pp[31][46] , \pp[31][45] , 
    \pp[31][44] , \pp[31][43] , \pp[31][42] , \pp[31][41] , \pp[31][40] , \pp[31][39] , 
    \pp[31][38] , \pp[31][37] , \pp[31][36] , \pp[31][35] , \pp[31][34] , \pp[31][33] , 
    \pp[31][32] , \pp[31][31] , uc_4227, uc_4228, uc_4229, uc_4230, uc_4231, uc_4232, 
    uc_4233, uc_4234, uc_4235, uc_4236, uc_4237, uc_4238, uc_4239, uc_4240, uc_4241, 
    uc_4242, uc_4243, uc_4244, uc_4245, uc_4246, uc_4247, uc_4248, uc_4249, uc_4250, 
    uc_4251, uc_4252, uc_4253, uc_4254, uc_4255, uc_4256, uc_4257}));
CSA__5_194 CSA16 (.u ({\sums[16][63] , \sums[16][62] , \sums[16][61] , \sums[16][60] , 
    \sums[16][59] , \sums[16][58] , \sums[16][57] , \sums[16][56] , \sums[16][55] , 
    \sums[16][54] , \sums[16][53] , \sums[16][52] , \sums[16][51] , \sums[16][50] , 
    \sums[16][49] , \sums[16][48] , \sums[16][47] , \sums[16][46] , \sums[16][45] , 
    \sums[16][44] , \sums[16][43] , \sums[16][42] , \sums[16][41] , \sums[16][40] , 
    \sums[16][39] , \sums[16][38] , \sums[16][37] , \sums[16][36] , \sums[16][35] , 
    \sums[16][34] , \sums[16][33] , \sums[16][32] , \sums[16][31] , \sums[16][30] , 
    \sums[16][29] , uc_4107, uc_4108, uc_4109, uc_4110, uc_4111, uc_4112, uc_4113, 
    uc_4114, uc_4115, uc_4116, uc_4117, uc_4118, uc_4119, uc_4120, uc_4121, uc_4122, 
    uc_4123, uc_4124, uc_4125, uc_4126, uc_4127, uc_4128, uc_4129, uc_4130, uc_4131, 
    uc_4132, uc_4133, uc_4134, uc_4135}), .v ({\couts[16][63] , \couts[16][62] , 
    \couts[16][61] , \couts[16][60] , \couts[16][59] , \couts[16][58] , \couts[16][57] , 
    \couts[16][56] , \couts[16][55] , \couts[16][54] , \couts[16][53] , \couts[16][52] , 
    \couts[16][51] , \couts[16][50] , \couts[16][49] , \couts[16][48] , \couts[16][47] , 
    \couts[16][46] , \couts[16][45] , \couts[16][44] , \couts[16][43] , \couts[16][42] , 
    \couts[16][41] , \couts[16][40] , \couts[16][39] , \couts[16][38] , \couts[16][37] , 
    \couts[16][36] , \couts[16][35] , \couts[16][34] , \couts[16][33] , \couts[16][32] , 
    \couts[16][31] , \couts[16][30] , uc_4136, uc_4137, uc_4138, uc_4139, uc_4140, 
    uc_4141, uc_4142, uc_4143, uc_4144, uc_4145, uc_4146, uc_4147, uc_4148, uc_4149, 
    uc_4150, uc_4151, uc_4152, uc_4153, uc_4154, uc_4155, uc_4156, uc_4157, uc_4158, 
    uc_4159, uc_4160, uc_4161, uc_4162, uc_4163, uc_4164, uc_4165}), .x ({\sums[9][63] , 
    \sums[9][62] , \sums[9][61] , \sums[9][60] , \sums[9][59] , \sums[9][58] , \sums[9][57] , 
    \sums[9][56] , \sums[9][55] , \sums[9][54] , \sums[9][53] , \sums[9][52] , \sums[9][51] , 
    \sums[9][50] , \sums[9][49] , \sums[9][48] , \sums[9][47] , \sums[9][46] , \sums[9][45] , 
    \sums[9][44] , \sums[9][43] , \sums[9][42] , \sums[9][41] , \sums[9][40] , \sums[9][39] , 
    \sums[9][38] , \sums[9][37] , \sums[9][36] , \sums[9][35] , \sums[9][34] , \sums[9][33] , 
    \sums[9][32] , \sums[9][31] , \sums[9][30] , \sums[9][29] , uc_4017, uc_4018, 
    uc_4019, uc_4020, uc_4021, uc_4022, uc_4023, uc_4024, uc_4025, uc_4026, uc_4027, 
    uc_4028, uc_4029, uc_4030, uc_4031, uc_4032, uc_4033, uc_4034, uc_4035, uc_4036, 
    uc_4037, uc_4038, uc_4039, uc_4040, uc_4041, uc_4042, uc_4043, uc_4044, uc_4045})
    , .y ({\couts[9][63] , \couts[9][62] , \couts[9][61] , \couts[9][60] , \couts[9][59] , 
    \couts[9][58] , \couts[9][57] , \couts[9][56] , \couts[9][55] , \couts[9][54] , 
    \couts[9][53] , \couts[9][52] , \couts[9][51] , \couts[9][50] , \couts[9][49] , 
    \couts[9][48] , \couts[9][47] , \couts[9][46] , \couts[9][45] , \couts[9][44] , 
    \couts[9][43] , \couts[9][42] , \couts[9][41] , \couts[9][40] , \couts[9][39] , 
    \couts[9][38] , \couts[9][37] , \couts[9][36] , \couts[9][35] , \couts[9][34] , 
    \couts[9][33] , \couts[9][32] , \couts[9][31] , \couts[9][30] , \couts[9][29] , 
    uc_4046, uc_4047, uc_4048, uc_4049, uc_4050, uc_4051, uc_4052, uc_4053, uc_4054, 
    uc_4055, uc_4056, uc_4057, uc_4058, uc_4059, uc_4060, uc_4061, uc_4062, uc_4063, 
    uc_4064, uc_4065, uc_4066, uc_4067, uc_4068, uc_4069, uc_4070, uc_4071, uc_4072, 
    uc_4073, uc_4074}), .z ({uc_4075, \pp[30][63] , uc_4076, \pp[30][60] , \pp[30][59] , 
    \pp[30][58] , \pp[30][57] , \pp[30][56] , \pp[30][55] , \pp[30][54] , \pp[30][53] , 
    \pp[30][52] , \pp[30][51] , \pp[30][50] , \pp[30][49] , \pp[30][48] , \pp[30][47] , 
    \pp[30][46] , \pp[30][45] , \pp[30][44] , \pp[30][43] , \pp[30][42] , \pp[30][41] , 
    \pp[30][40] , \pp[30][39] , \pp[30][38] , \pp[30][37] , \pp[30][36] , \pp[30][35] , 
    \pp[30][34] , \pp[30][33] , \pp[30][32] , \pp[30][31] , \pp[30][30] , uc_4077, 
    uc_4078, uc_4079, uc_4080, uc_4081, uc_4082, uc_4083, uc_4084, uc_4085, uc_4086, 
    uc_4087, uc_4088, uc_4089, uc_4090, uc_4091, uc_4092, uc_4093, uc_4094, uc_4095, 
    uc_4096, uc_4097, uc_4098, uc_4099, uc_4100, uc_4101, uc_4102, uc_4103, uc_4104, 
    uc_4105, uc_4106}));
CSA__5_191 CSA9 (.u ({\sums[9][63] , \sums[9][62] , \sums[9][61] , \sums[9][60] , 
    \sums[9][59] , \sums[9][58] , \sums[9][57] , \sums[9][56] , \sums[9][55] , \sums[9][54] , 
    \sums[9][53] , \sums[9][52] , \sums[9][51] , \sums[9][50] , \sums[9][49] , \sums[9][48] , 
    \sums[9][47] , \sums[9][46] , \sums[9][45] , \sums[9][44] , \sums[9][43] , \sums[9][42] , 
    \sums[9][41] , \sums[9][40] , \sums[9][39] , \sums[9][38] , \sums[9][37] , \sums[9][36] , 
    \sums[9][35] , \sums[9][34] , \sums[9][33] , \sums[9][32] , \sums[9][31] , \sums[9][30] , 
    \sums[9][29] , \sums[9][28] , uc_3960, uc_3961, uc_3962, uc_3963, uc_3964, uc_3965, 
    uc_3966, uc_3967, uc_3968, uc_3969, uc_3970, uc_3971, uc_3972, uc_3973, uc_3974, 
    uc_3975, uc_3976, uc_3977, uc_3978, uc_3979, uc_3980, uc_3981, uc_3982, uc_3983, 
    uc_3984, uc_3985, uc_3986, uc_3987}), .v ({\couts[9][63] , \couts[9][62] , \couts[9][61] , 
    \couts[9][60] , \couts[9][59] , \couts[9][58] , \couts[9][57] , \couts[9][56] , 
    \couts[9][55] , \couts[9][54] , \couts[9][53] , \couts[9][52] , \couts[9][51] , 
    \couts[9][50] , \couts[9][49] , \couts[9][48] , \couts[9][47] , \couts[9][46] , 
    \couts[9][45] , \couts[9][44] , \couts[9][43] , \couts[9][42] , \couts[9][41] , 
    \couts[9][40] , \couts[9][39] , \couts[9][38] , \couts[9][37] , \couts[9][36] , 
    \couts[9][35] , \couts[9][34] , \couts[9][33] , \couts[9][32] , \couts[9][31] , 
    \couts[9][30] , \couts[9][29] , uc_3988, uc_3989, uc_3990, uc_3991, uc_3992, 
    uc_3993, uc_3994, uc_3995, uc_3996, uc_3997, uc_3998, uc_3999, uc_4000, uc_4001, 
    uc_4002, uc_4003, uc_4004, uc_4005, uc_4006, uc_4007, uc_4008, uc_4009, uc_4010, 
    uc_4011, uc_4012, uc_4013, uc_4014, uc_4015, uc_4016}), .x ({\pp[27][58] , \pp[27][58] , 
    \pp[27][58] , \pp[27][58] , \pp[27][58] , \pp[27][58] , \pp[27][57] , \pp[27][56] , 
    \pp[27][55] , \pp[27][54] , \pp[27][53] , \pp[27][52] , \pp[27][51] , \pp[27][50] , 
    \pp[27][49] , \pp[27][48] , \pp[27][47] , \pp[27][46] , \pp[27][45] , \pp[27][44] , 
    \pp[27][43] , \pp[27][42] , \pp[27][41] , \pp[27][40] , \pp[27][39] , \pp[27][38] , 
    \pp[27][37] , \pp[27][36] , \pp[27][35] , \pp[27][34] , \pp[27][33] , \pp[27][32] , 
    \pp[27][31] , \pp[27][30] , \pp[27][29] , \pp[27][28] , uc_3868, uc_3869, uc_3870, 
    uc_3871, uc_3872, uc_3873, uc_3874, uc_3875, uc_3876, uc_3877, uc_3878, uc_3879, 
    uc_3880, uc_3881, uc_3882, uc_3883, uc_3884, uc_3885, uc_3886, uc_3887, uc_3888, 
    uc_3889, uc_3890, uc_3891, uc_3892, uc_3893, uc_3894, uc_3895}), .y ({uc_3896, 
    \pp[28][63] , uc_3897, uc_3898, uc_3899, \pp[28][58] , \pp[28][57] , \pp[28][56] , 
    \pp[28][55] , \pp[28][54] , \pp[28][53] , \pp[28][52] , \pp[28][51] , \pp[28][50] , 
    \pp[28][49] , \pp[28][48] , \pp[28][47] , \pp[28][46] , \pp[28][45] , \pp[28][44] , 
    \pp[28][43] , \pp[28][42] , \pp[28][41] , \pp[28][40] , \pp[28][39] , \pp[28][38] , 
    \pp[28][37] , \pp[28][36] , \pp[28][35] , \pp[28][34] , \pp[28][33] , \pp[28][32] , 
    \pp[28][31] , \pp[28][30] , \pp[28][29] , \pp[28][28] , uc_3900, uc_3901, uc_3902, 
    uc_3903, uc_3904, uc_3905, uc_3906, uc_3907, uc_3908, uc_3909, uc_3910, uc_3911, 
    uc_3912, uc_3913, uc_3914, uc_3915, uc_3916, uc_3917, uc_3918, uc_3919, uc_3920, 
    uc_3921, uc_3922, uc_3923, uc_3924, uc_3925, uc_3926, uc_3927}), .z ({uc_3928, 
    \pp[29][63] , uc_3929, uc_3930, \pp[29][59] , \pp[29][58] , \pp[29][57] , \pp[29][56] , 
    \pp[29][55] , \pp[29][54] , \pp[29][53] , \pp[29][52] , \pp[29][51] , \pp[29][50] , 
    \pp[29][49] , \pp[29][48] , \pp[29][47] , \pp[29][46] , \pp[29][45] , \pp[29][44] , 
    \pp[29][43] , \pp[29][42] , \pp[29][41] , \pp[29][40] , \pp[29][39] , \pp[29][38] , 
    \pp[29][37] , \pp[29][36] , \pp[29][35] , \pp[29][34] , \pp[29][33] , \pp[29][32] , 
    \pp[29][31] , \pp[29][30] , \pp[29][29] , uc_3931, uc_3932, uc_3933, uc_3934, 
    uc_3935, uc_3936, uc_3937, uc_3938, uc_3939, uc_3940, uc_3941, uc_3942, uc_3943, 
    uc_3944, uc_3945, uc_3946, uc_3947, uc_3948, uc_3949, uc_3950, uc_3951, uc_3952, 
    uc_3953, uc_3954, uc_3955, uc_3956, uc_3957, uc_3958, uc_3959}));
CSA__0_78 CSA20 (.u ({\sums[20][59] , uc_3814, uc_3815, uc_3816, uc_3817, \sums[20][58] , 
    \sums[20][57] , \sums[20][56] , \sums[20][55] , \sums[20][54] , \sums[20][53] , 
    \sums[20][52] , \sums[20][51] , \sums[20][50] , \sums[20][49] , \sums[20][48] , 
    \sums[20][47] , \sums[20][46] , \sums[20][45] , \sums[20][44] , \sums[20][43] , 
    \sums[20][42] , \sums[20][41] , \sums[20][40] , \sums[20][39] , \sums[20][38] , 
    \sums[20][37] , \sums[20][36] , \sums[20][35] , \sums[20][34] , \sums[20][33] , 
    \sums[20][32] , \sums[20][31] , \sums[20][30] , \sums[20][29] , \sums[20][28] , 
    \sums[20][27] , \sums[20][26] , \sums[20][25] , \sums[20][24] , \sums[20][23] , 
    uc_3818, uc_3819, uc_3820, uc_3821, uc_3822, uc_3823, uc_3824, uc_3825, uc_3826, 
    uc_3827, uc_3828, uc_3829, uc_3830, uc_3831, uc_3832, uc_3833, uc_3834, uc_3835, 
    uc_3836, uc_3837, uc_3838, uc_3839, uc_3840}), .v ({\couts[20][63] , uc_3841, 
    uc_3842, uc_3843, \couts[20][59] , \couts[20][58] , \couts[20][57] , \couts[20][56] , 
    \couts[20][55] , \couts[20][54] , \couts[20][53] , \couts[20][52] , \couts[20][51] , 
    \couts[20][50] , \couts[20][49] , \couts[20][48] , \couts[20][47] , \couts[20][46] , 
    \couts[20][45] , \couts[20][44] , \couts[20][43] , \couts[20][42] , \couts[20][41] , 
    \couts[20][40] , \couts[20][39] , \couts[20][38] , \couts[20][37] , \couts[20][36] , 
    \couts[20][35] , \couts[20][34] , \couts[20][33] , \couts[20][32] , \couts[20][31] , 
    \couts[20][30] , \couts[20][29] , \couts[20][28] , \couts[20][27] , \couts[20][26] , 
    \couts[20][25] , \couts[20][24] , uc_3844, uc_3845, uc_3846, uc_3847, uc_3848, 
    uc_3849, uc_3850, uc_3851, uc_3852, uc_3853, uc_3854, uc_3855, uc_3856, uc_3857, 
    uc_3858, uc_3859, uc_3860, uc_3861, uc_3862, uc_3863, uc_3864, uc_3865, uc_3866, 
    uc_3867}), .x ({\couts[14][63] , uc_3726, uc_3727, uc_3728, uc_3729, uc_3730, 
    uc_3731, uc_3732, uc_3733, \couts[14][54] , \couts[14][53] , \couts[14][52] , 
    \couts[14][51] , \couts[14][50] , \couts[14][49] , \couts[14][48] , \couts[14][47] , 
    \couts[14][46] , \couts[14][45] , \couts[14][44] , \couts[14][43] , \couts[14][42] , 
    \couts[14][41] , \couts[14][40] , \couts[14][39] , \couts[14][38] , \couts[14][37] , 
    \couts[14][36] , \couts[14][35] , \couts[14][34] , \couts[14][33] , \couts[14][32] , 
    \couts[14][31] , \couts[14][30] , \couts[14][29] , \couts[14][28] , \couts[14][27] , 
    \couts[14][26] , \couts[14][25] , \couts[14][24] , \couts[14][23] , uc_3734, 
    uc_3735, uc_3736, uc_3737, uc_3738, uc_3739, uc_3740, uc_3741, uc_3742, uc_3743, 
    uc_3744, uc_3745, uc_3746, uc_3747, uc_3748, uc_3749, uc_3750, uc_3751, uc_3752, 
    uc_3753, uc_3754, uc_3755, uc_3756}), .y ({\sums[15][63] , uc_3757, uc_3758, 
    uc_3759, uc_3760, uc_3761, \sums[15][57] , \sums[15][56] , \sums[15][55] , \sums[15][54] , 
    \sums[15][53] , \sums[15][52] , \sums[15][51] , \sums[15][50] , \sums[15][49] , 
    \sums[15][48] , \sums[15][47] , \sums[15][46] , \sums[15][45] , \sums[15][44] , 
    \sums[15][43] , \sums[15][42] , \sums[15][41] , \sums[15][40] , \sums[15][39] , 
    \sums[15][38] , \sums[15][37] , \sums[15][36] , \sums[15][35] , \sums[15][34] , 
    \sums[15][33] , \sums[15][32] , \sums[15][31] , \sums[15][30] , \sums[15][29] , 
    \sums[15][28] , \sums[15][27] , \sums[15][26] , \sums[15][25] , \sums[15][24] , 
    \couts[7][23] , uc_3762, uc_3763, uc_3764, uc_3765, uc_3766, uc_3767, uc_3768, 
    uc_3769, uc_3770, uc_3771, uc_3772, uc_3773, uc_3774, uc_3775, uc_3776, uc_3777, 
    uc_3778, uc_3779, uc_3780, uc_3781, uc_3782, uc_3783, uc_3784}), .z ({\couts[15][63] , 
    uc_3785, uc_3786, uc_3787, uc_3788, \couts[15][58] , \couts[15][57] , \couts[15][56] , 
    \couts[15][55] , \couts[15][54] , \couts[15][53] , \couts[15][52] , \couts[15][51] , 
    \couts[15][50] , \couts[15][49] , \couts[15][48] , \couts[15][47] , \couts[15][46] , 
    \couts[15][45] , \couts[15][44] , \couts[15][43] , \couts[15][42] , \couts[15][41] , 
    \couts[15][40] , \couts[15][39] , \couts[15][38] , \couts[15][37] , \couts[15][36] , 
    \couts[15][35] , \couts[15][34] , \couts[15][33] , \couts[15][32] , \couts[15][31] , 
    \couts[15][30] , \couts[15][29] , \couts[15][28] , \couts[15][27] , \couts[15][26] , 
    \couts[15][25] , uc_3789, uc_3790, uc_3791, uc_3792, uc_3793, uc_3794, uc_3795, 
    uc_3796, uc_3797, uc_3798, uc_3799, uc_3800, uc_3801, uc_3802, uc_3803, uc_3804, 
    uc_3805, uc_3806, uc_3807, uc_3808, uc_3809, uc_3810, uc_3811, uc_3812, uc_3813}));
CSA__4_20 CSA15 (.u ({\sums[15][63] , uc_3668, uc_3669, uc_3670, uc_3671, uc_3672, 
    \sums[15][57] , \sums[15][56] , \sums[15][55] , \sums[15][54] , \sums[15][53] , 
    \sums[15][52] , \sums[15][51] , \sums[15][50] , \sums[15][49] , \sums[15][48] , 
    \sums[15][47] , \sums[15][46] , \sums[15][45] , \sums[15][44] , \sums[15][43] , 
    \sums[15][42] , \sums[15][41] , \sums[15][40] , \sums[15][39] , \sums[15][38] , 
    \sums[15][37] , \sums[15][36] , \sums[15][35] , \sums[15][34] , \sums[15][33] , 
    \sums[15][32] , \sums[15][31] , \sums[15][30] , \sums[15][29] , \sums[15][28] , 
    \sums[15][27] , \sums[15][26] , \sums[15][25] , \sums[15][24] , uc_3673, uc_3674, 
    uc_3675, uc_3676, uc_3677, uc_3678, uc_3679, uc_3680, uc_3681, uc_3682, uc_3683, 
    uc_3684, uc_3685, uc_3686, uc_3687, uc_3688, uc_3689, uc_3690, uc_3691, uc_3692, 
    uc_3693, uc_3694, uc_3695, uc_3696}), .v ({\couts[15][63] , uc_3697, uc_3698, 
    uc_3699, uc_3700, \couts[15][58] , \couts[15][57] , \couts[15][56] , \couts[15][55] , 
    \couts[15][54] , \couts[15][53] , \couts[15][52] , \couts[15][51] , \couts[15][50] , 
    \couts[15][49] , \couts[15][48] , \couts[15][47] , \couts[15][46] , \couts[15][45] , 
    \couts[15][44] , \couts[15][43] , \couts[15][42] , \couts[15][41] , \couts[15][40] , 
    \couts[15][39] , \couts[15][38] , \couts[15][37] , \couts[15][36] , \couts[15][35] , 
    \couts[15][34] , \couts[15][33] , \couts[15][32] , \couts[15][31] , \couts[15][30] , 
    \couts[15][29] , \couts[15][28] , \couts[15][27] , \couts[15][26] , \couts[15][25] , 
    uc_3701, uc_3702, uc_3703, uc_3704, uc_3705, uc_3706, uc_3707, uc_3708, uc_3709, 
    uc_3710, uc_3711, uc_3712, uc_3713, uc_3714, uc_3715, uc_3716, uc_3717, uc_3718, 
    uc_3719, uc_3720, uc_3721, uc_3722, uc_3723, uc_3724, uc_3725}), .x ({\couts[7][63] , 
    uc_3575, uc_3576, uc_3577, uc_3578, uc_3579, uc_3580, uc_3581, uc_3582, \couts[7][54] , 
    \couts[7][53] , \couts[7][52] , \couts[7][51] , \couts[7][50] , \couts[7][49] , 
    \couts[7][48] , \couts[7][47] , \couts[7][46] , \couts[7][45] , \couts[7][44] , 
    \couts[7][43] , \couts[7][42] , \couts[7][41] , \couts[7][40] , \couts[7][39] , 
    \couts[7][38] , \couts[7][37] , \couts[7][36] , \couts[7][35] , \couts[7][34] , 
    \couts[7][33] , \couts[7][32] , \couts[7][31] , \couts[7][30] , \couts[7][29] , 
    \couts[7][28] , \couts[7][27] , \couts[7][26] , \couts[7][25] , \couts[7][24] , 
    uc_3583, uc_3584, uc_3585, uc_3586, uc_3587, uc_3588, uc_3589, uc_3590, uc_3591, 
    uc_3592, uc_3593, uc_3594, uc_3595, uc_3596, uc_3597, uc_3598, uc_3599, uc_3600, 
    uc_3601, uc_3602, uc_3603, uc_3604, uc_3605, uc_3606}), .y ({\sums[8][63] , uc_3607, 
    uc_3608, uc_3609, uc_3610, uc_3611, uc_3612, \sums[8][56] , \sums[8][55] , \sums[8][54] , 
    \sums[8][53] , \sums[8][52] , \sums[8][51] , \sums[8][50] , \sums[8][49] , \sums[8][48] , 
    \sums[8][47] , \sums[8][46] , \sums[8][45] , \sums[8][44] , \sums[8][43] , \sums[8][42] , 
    \sums[8][41] , \sums[8][40] , \sums[8][39] , \sums[8][38] , \sums[8][37] , \sums[8][36] , 
    \sums[8][35] , \sums[8][34] , \sums[8][33] , \sums[8][32] , \sums[8][31] , \sums[8][30] , 
    \sums[8][29] , \sums[8][28] , \sums[8][27] , \sums[8][26] , \sums[8][25] , \pp[24][24] , 
    uc_3613, uc_3614, uc_3615, uc_3616, uc_3617, uc_3618, uc_3619, uc_3620, uc_3621, 
    uc_3622, uc_3623, uc_3624, uc_3625, uc_3626, uc_3627, uc_3628, uc_3629, uc_3630, 
    uc_3631, uc_3632, uc_3633, uc_3634, uc_3635, uc_3636}), .z ({\couts[8][63] , 
    uc_3637, uc_3638, uc_3639, uc_3640, uc_3641, \couts[8][57] , \couts[8][56] , 
    \couts[8][55] , \couts[8][54] , \couts[8][53] , \couts[8][52] , \couts[8][51] , 
    \couts[8][50] , \couts[8][49] , \couts[8][48] , \couts[8][47] , \couts[8][46] , 
    \couts[8][45] , \couts[8][44] , \couts[8][43] , \couts[8][42] , \couts[8][41] , 
    \couts[8][40] , \couts[8][39] , \couts[8][38] , \couts[8][37] , \couts[8][36] , 
    \couts[8][35] , \couts[8][34] , \couts[8][33] , \couts[8][32] , \couts[8][31] , 
    \couts[8][30] , \couts[8][29] , \couts[8][28] , \couts[8][27] , \couts[8][26] , 
    uc_3642, uc_3643, uc_3644, uc_3645, uc_3646, uc_3647, uc_3648, uc_3649, uc_3650, 
    uc_3651, uc_3652, uc_3653, uc_3654, uc_3655, uc_3656, uc_3657, uc_3658, uc_3659, 
    uc_3660, uc_3661, uc_3662, uc_3663, uc_3664, uc_3665, uc_3666, uc_3667}));
CSA__4_17 CSA8 (.u ({\sums[8][63] , uc_3513, uc_3514, uc_3515, uc_3516, uc_3517, 
    uc_3518, \sums[8][56] , \sums[8][55] , \sums[8][54] , \sums[8][53] , \sums[8][52] , 
    \sums[8][51] , \sums[8][50] , \sums[8][49] , \sums[8][48] , \sums[8][47] , \sums[8][46] , 
    \sums[8][45] , \sums[8][44] , \sums[8][43] , \sums[8][42] , \sums[8][41] , \sums[8][40] , 
    \sums[8][39] , \sums[8][38] , \sums[8][37] , \sums[8][36] , \sums[8][35] , \sums[8][34] , 
    \sums[8][33] , \sums[8][32] , \sums[8][31] , \sums[8][30] , \sums[8][29] , \sums[8][28] , 
    \sums[8][27] , \sums[8][26] , \sums[8][25] , uc_3519, uc_3520, uc_3521, uc_3522, 
    uc_3523, uc_3524, uc_3525, uc_3526, uc_3527, uc_3528, uc_3529, uc_3530, uc_3531, 
    uc_3532, uc_3533, uc_3534, uc_3535, uc_3536, uc_3537, uc_3538, uc_3539, uc_3540, 
    uc_3541, uc_3542, uc_3543}), .v ({\couts[8][63] , uc_3544, uc_3545, uc_3546, 
    uc_3547, uc_3548, \couts[8][57] , \couts[8][56] , \couts[8][55] , \couts[8][54] , 
    \couts[8][53] , \couts[8][52] , \couts[8][51] , \couts[8][50] , \couts[8][49] , 
    \couts[8][48] , \couts[8][47] , \couts[8][46] , \couts[8][45] , \couts[8][44] , 
    \couts[8][43] , \couts[8][42] , \couts[8][41] , \couts[8][40] , \couts[8][39] , 
    \couts[8][38] , \couts[8][37] , \couts[8][36] , \couts[8][35] , \couts[8][34] , 
    \couts[8][33] , \couts[8][32] , \couts[8][31] , \couts[8][30] , \couts[8][29] , 
    \couts[8][28] , \couts[8][27] , \couts[8][26] , uc_3549, uc_3550, uc_3551, uc_3552, 
    uc_3553, uc_3554, uc_3555, uc_3556, uc_3557, uc_3558, uc_3559, uc_3560, uc_3561, 
    uc_3562, uc_3563, uc_3564, uc_3565, uc_3566, uc_3567, uc_3568, uc_3569, uc_3570, 
    uc_3571, uc_3572, uc_3573, uc_3574}), .x ({\pp[24][63] , uc_3416, uc_3417, uc_3418, 
    uc_3419, uc_3420, uc_3421, uc_3422, uc_3423, \pp[24][54] , \pp[24][53] , \pp[24][52] , 
    \pp[24][51] , \pp[24][50] , \pp[24][49] , \pp[24][48] , \pp[24][47] , \pp[24][46] , 
    \pp[24][45] , \pp[24][44] , \pp[24][43] , \pp[24][42] , \pp[24][41] , \pp[24][40] , 
    \pp[24][39] , \pp[24][38] , \pp[24][37] , \pp[24][36] , \pp[24][35] , \pp[24][34] , 
    \pp[24][33] , \pp[24][32] , \pp[24][31] , \pp[24][30] , \pp[24][29] , \pp[24][28] , 
    \pp[24][27] , \pp[24][26] , \pp[24][25] , uc_3424, uc_3425, uc_3426, uc_3427, 
    uc_3428, uc_3429, uc_3430, uc_3431, uc_3432, uc_3433, uc_3434, uc_3435, uc_3436, 
    uc_3437, uc_3438, uc_3439, uc_3440, uc_3441, uc_3442, uc_3443, uc_3444, uc_3445, 
    uc_3446, uc_3447, uc_3448}), .y ({\pp[25][63] , uc_3449, uc_3450, uc_3451, uc_3452, 
    uc_3453, uc_3454, uc_3455, \pp[25][55] , \pp[25][54] , \pp[25][53] , \pp[25][52] , 
    \pp[25][51] , \pp[25][50] , \pp[25][49] , \pp[25][48] , \pp[25][47] , \pp[25][46] , 
    \pp[25][45] , \pp[25][44] , \pp[25][43] , \pp[25][42] , \pp[25][41] , \pp[25][40] , 
    \pp[25][39] , \pp[25][38] , \pp[25][37] , \pp[25][36] , \pp[25][35] , \pp[25][34] , 
    \pp[25][33] , \pp[25][32] , \pp[25][31] , \pp[25][30] , \pp[25][29] , \pp[25][28] , 
    \pp[25][27] , \pp[25][26] , \pp[25][25] , uc_3456, uc_3457, uc_3458, uc_3459, 
    uc_3460, uc_3461, uc_3462, uc_3463, uc_3464, uc_3465, uc_3466, uc_3467, uc_3468, 
    uc_3469, uc_3470, uc_3471, uc_3472, uc_3473, uc_3474, uc_3475, uc_3476, uc_3477, 
    uc_3478, uc_3479, uc_3480}), .z ({\pp[26][63] , uc_3481, uc_3482, uc_3483, uc_3484, 
    uc_3485, uc_3486, \pp[26][56] , \pp[26][55] , \pp[26][54] , \pp[26][53] , \pp[26][52] , 
    \pp[26][51] , \pp[26][50] , \pp[26][49] , \pp[26][48] , \pp[26][47] , \pp[26][46] , 
    \pp[26][45] , \pp[26][44] , \pp[26][43] , \pp[26][42] , \pp[26][41] , \pp[26][40] , 
    \pp[26][39] , \pp[26][38] , \pp[26][37] , \pp[26][36] , \pp[26][35] , \pp[26][34] , 
    \pp[26][33] , \pp[26][32] , \pp[26][31] , \pp[26][30] , \pp[26][29] , \pp[26][28] , 
    \pp[26][27] , \pp[26][26] , uc_3487, uc_3488, uc_3489, uc_3490, uc_3491, uc_3492, 
    uc_3493, uc_3494, uc_3495, uc_3496, uc_3497, uc_3498, uc_3499, uc_3500, uc_3501, 
    uc_3502, uc_3503, uc_3504, uc_3505, uc_3506, uc_3507, uc_3508, uc_3509, uc_3510, 
    uc_3511, uc_3512}));
CSA__4_14 CSA6 (.u ({\sums[6][63] , uc_3354, uc_3355, uc_3356, uc_3357, uc_3358, 
    uc_3359, uc_3360, uc_3361, uc_3362, uc_3363, uc_3364, uc_3365, \sums[6][50] , 
    \sums[6][49] , \sums[6][48] , \sums[6][47] , \sums[6][46] , \sums[6][45] , \sums[6][44] , 
    \sums[6][43] , \sums[6][42] , \sums[6][41] , \sums[6][40] , \sums[6][39] , \sums[6][38] , 
    \sums[6][37] , \sums[6][36] , \sums[6][35] , \sums[6][34] , \sums[6][33] , \sums[6][32] , 
    \sums[6][31] , \sums[6][30] , \sums[6][29] , \sums[6][28] , \sums[6][27] , \sums[6][26] , 
    \sums[6][25] , \sums[6][24] , \sums[6][23] , \sums[6][22] , \sums[6][21] , \sums[6][20] , 
    \sums[6][19] , uc_3366, uc_3367, uc_3368, uc_3369, uc_3370, uc_3371, uc_3372, 
    uc_3373, uc_3374, uc_3375, uc_3376, uc_3377, uc_3378, uc_3379, uc_3380, uc_3381, 
    uc_3382, uc_3383, uc_3384}), .v ({\couts[6][63] , uc_3385, uc_3386, uc_3387, 
    uc_3388, uc_3389, uc_3390, uc_3391, uc_3392, uc_3393, uc_3394, uc_3395, \couts[6][51] , 
    \couts[6][50] , \couts[6][49] , \couts[6][48] , \couts[6][47] , \couts[6][46] , 
    \couts[6][45] , \couts[6][44] , \couts[6][43] , \couts[6][42] , \couts[6][41] , 
    \couts[6][40] , \couts[6][39] , \couts[6][38] , \couts[6][37] , \couts[6][36] , 
    \couts[6][35] , \couts[6][34] , \couts[6][33] , \couts[6][32] , \couts[6][31] , 
    \couts[6][30] , \couts[6][29] , \couts[6][28] , \couts[6][27] , \couts[6][26] , 
    \couts[6][25] , \couts[6][24] , \couts[6][23] , \couts[6][22] , \couts[6][21] , 
    \couts[6][20] , uc_3396, uc_3397, uc_3398, uc_3399, uc_3400, uc_3401, uc_3402, 
    uc_3403, uc_3404, uc_3405, uc_3406, uc_3407, uc_3408, uc_3409, uc_3410, uc_3411, 
    uc_3412, uc_3413, uc_3414, uc_3415}), .x ({uc_3257, \pp[18][63] , uc_3258, uc_3259, 
    uc_3260, uc_3261, uc_3262, uc_3263, uc_3264, uc_3265, uc_3266, uc_3267, uc_3268, 
    uc_3269, uc_3270, \pp[18][48] , \pp[18][47] , \pp[18][46] , \pp[18][45] , \pp[18][44] , 
    \pp[18][43] , \pp[18][42] , \pp[18][41] , \pp[18][40] , \pp[18][39] , \pp[18][38] , 
    \pp[18][37] , \pp[18][36] , \pp[18][35] , \pp[18][34] , \pp[18][33] , \pp[18][32] , 
    \pp[18][31] , \pp[18][30] , \pp[18][29] , \pp[18][28] , \pp[18][27] , \pp[18][26] , 
    \pp[18][25] , \pp[18][24] , \pp[18][23] , \pp[18][22] , \pp[18][21] , \pp[18][20] , 
    \pp[18][19] , uc_3271, uc_3272, uc_3273, uc_3274, uc_3275, uc_3276, uc_3277, 
    uc_3278, uc_3279, uc_3280, uc_3281, uc_3282, uc_3283, uc_3284, uc_3285, uc_3286, 
    uc_3287, uc_3288, uc_3289}), .y ({uc_3290, \pp[19][63] , uc_3291, uc_3292, uc_3293, 
    uc_3294, uc_3295, uc_3296, uc_3297, uc_3298, uc_3299, uc_3300, uc_3301, uc_3302, 
    \pp[19][49] , \pp[19][48] , \pp[19][47] , \pp[19][46] , \pp[19][45] , \pp[19][44] , 
    \pp[19][43] , \pp[19][42] , \pp[19][41] , \pp[19][40] , \pp[19][39] , \pp[19][38] , 
    \pp[19][37] , \pp[19][36] , \pp[19][35] , \pp[19][34] , \pp[19][33] , \pp[19][32] , 
    \pp[19][31] , \pp[19][30] , \pp[19][29] , \pp[19][28] , \pp[19][27] , \pp[19][26] , 
    \pp[19][25] , \pp[19][24] , \pp[19][23] , \pp[19][22] , \pp[19][21] , \pp[19][20] , 
    \pp[19][19] , uc_3303, uc_3304, uc_3305, uc_3306, uc_3307, uc_3308, uc_3309, 
    uc_3310, uc_3311, uc_3312, uc_3313, uc_3314, uc_3315, uc_3316, uc_3317, uc_3318, 
    uc_3319, uc_3320, uc_3321}), .z ({uc_3322, \pp[20][63] , uc_3323, uc_3324, uc_3325, 
    uc_3326, uc_3327, uc_3328, uc_3329, uc_3330, uc_3331, uc_3332, uc_3333, \pp[20][50] , 
    \pp[20][49] , \pp[20][48] , \pp[20][47] , \pp[20][46] , \pp[20][45] , \pp[20][44] , 
    \pp[20][43] , \pp[20][42] , \pp[20][41] , \pp[20][40] , \pp[20][39] , \pp[20][38] , 
    \pp[20][37] , \pp[20][36] , \pp[20][35] , \pp[20][34] , \pp[20][33] , \pp[20][32] , 
    \pp[20][31] , \pp[20][30] , \pp[20][29] , \pp[20][28] , \pp[20][27] , \pp[20][26] , 
    \pp[20][25] , \pp[20][24] , \pp[20][23] , \pp[20][22] , \pp[20][21] , \pp[20][20] , 
    uc_3334, uc_3335, uc_3336, uc_3337, uc_3338, uc_3339, uc_3340, uc_3341, uc_3342, 
    uc_3343, uc_3344, uc_3345, uc_3346, uc_3347, uc_3348, uc_3349, uc_3350, uc_3351, 
    uc_3352, uc_3353}));
CSA__4_11 CSA23 (.u ({\sums[23][63] , \sums[23][62] , \sums[23][61] , \sums[23][60] , 
    \sums[23][59] , \sums[23][58] , \sums[23][57] , \sums[23][56] , \sums[23][55] , 
    \sums[23][54] , \sums[23][53] , \sums[23][52] , \sums[23][51] , \sums[23][50] , 
    \sums[23][49] , \sums[23][48] , \sums[23][47] , \sums[23][46] , \sums[23][45] , 
    \sums[23][44] , \sums[23][43] , \sums[23][42] , \sums[23][41] , \sums[23][40] , 
    \sums[23][39] , \sums[23][38] , \sums[23][37] , \sums[23][36] , \sums[23][35] , 
    \sums[23][34] , \sums[23][33] , \sums[23][32] , \sums[23][31] , \sums[23][30] , 
    \sums[23][29] , \sums[23][28] , \sums[23][27] , \sums[23][26] , \sums[23][25] , 
    \sums[23][24] , \sums[23][23] , \sums[23][22] , \sums[23][21] , \sums[23][20] , 
    \sums[23][19] , \sums[23][18] , \sums[23][17] , \sums[23][16] , \sums[23][15] , 
    \sums[23][14] , uc_3228, uc_3229, uc_3230, uc_3231, uc_3232, uc_3233, uc_3234, 
    uc_3235, uc_3236, uc_3237, uc_3238, uc_3239, uc_3240, uc_3241}), .v ({\couts[23][63] , 
    \couts[23][62] , \couts[23][61] , \couts[23][60] , \couts[23][59] , \couts[23][58] , 
    \couts[23][57] , \couts[23][56] , \couts[23][55] , \couts[23][54] , \couts[23][53] , 
    \couts[23][52] , \couts[23][51] , \couts[23][50] , \couts[23][49] , \couts[23][48] , 
    \couts[23][47] , \couts[23][46] , \couts[23][45] , \couts[23][44] , \couts[23][43] , 
    \couts[23][42] , \couts[23][41] , \couts[23][40] , \couts[23][39] , \couts[23][38] , 
    \couts[23][37] , \couts[23][36] , \couts[23][35] , \couts[23][34] , \couts[23][33] , 
    \couts[23][32] , \couts[23][31] , \couts[23][30] , \couts[23][29] , \couts[23][28] , 
    \couts[23][27] , \couts[23][26] , \couts[23][25] , \couts[23][24] , \couts[23][23] , 
    \couts[23][22] , \couts[23][21] , \couts[23][20] , \couts[23][19] , \couts[23][18] , 
    \couts[23][17] , \couts[23][16] , \couts[23][15] , uc_3242, uc_3243, uc_3244, 
    uc_3245, uc_3246, uc_3247, uc_3248, uc_3249, uc_3250, uc_3251, uc_3252, uc_3253, 
    uc_3254, uc_3255, uc_3256}), .x ({\couts[18][63] , \couts[18][62] , \couts[18][61] , 
    \couts[18][60] , \couts[18][59] , \couts[18][58] , \couts[18][57] , \couts[18][56] , 
    \couts[18][55] , \couts[18][54] , \couts[18][53] , \couts[18][52] , \couts[18][51] , 
    \couts[18][50] , \couts[18][49] , \couts[18][48] , \couts[18][47] , \couts[18][46] , 
    \couts[18][45] , \couts[18][44] , \couts[18][43] , \couts[18][42] , \couts[18][41] , 
    \couts[18][40] , \couts[18][39] , \couts[18][38] , \couts[18][37] , \couts[18][36] , 
    \couts[18][35] , \couts[18][34] , \couts[18][33] , \couts[18][32] , \couts[18][31] , 
    \couts[18][30] , \couts[18][29] , \couts[18][28] , \couts[18][27] , \couts[18][26] , 
    \couts[18][25] , \couts[18][24] , \couts[18][23] , \couts[18][22] , \couts[18][21] , 
    \couts[18][20] , \couts[18][19] , \couts[18][18] , \couts[18][17] , \couts[18][16] , 
    \couts[18][15] , \couts[18][14] , uc_3166, uc_3167, uc_3168, uc_3169, uc_3170, 
    uc_3171, uc_3172, uc_3173, uc_3174, uc_3175, uc_3176, uc_3177, uc_3178, uc_3179})
    , .y ({\sums[19][63] , uc_3180, uc_3181, uc_3182, uc_3183, uc_3184, uc_3185, 
    uc_3186, uc_3187, uc_3188, \sums[19][53] , \sums[19][52] , \sums[19][51] , \sums[19][50] , 
    \sums[19][49] , \sums[19][48] , \sums[19][47] , \sums[19][46] , \sums[19][45] , 
    \sums[19][44] , \sums[19][43] , \sums[19][42] , \sums[19][41] , \sums[19][40] , 
    \sums[19][39] , \sums[19][38] , \sums[19][37] , \sums[19][36] , \sums[19][35] , 
    \sums[19][34] , \sums[19][33] , \sums[19][32] , \sums[19][31] , \sums[19][30] , 
    \sums[19][29] , \sums[19][28] , \sums[19][27] , \sums[19][26] , \sums[19][25] , 
    \sums[19][24] , \sums[19][23] , \sums[19][22] , \sums[19][21] , \sums[19][20] , 
    \sums[19][19] , \sums[19][18] , \sums[19][17] , \sums[19][16] , \sums[13][15] , 
    \sums[13][14] , uc_3189, uc_3190, uc_3191, uc_3192, uc_3193, uc_3194, uc_3195, 
    uc_3196, uc_3197, uc_3198, uc_3199, uc_3200, uc_3201, uc_3202}), .z ({\couts[19][63] , 
    uc_3203, uc_3204, uc_3205, uc_3206, uc_3207, uc_3208, uc_3209, uc_3210, \couts[19][54] , 
    \couts[19][53] , \couts[19][52] , \couts[19][51] , \couts[19][50] , \couts[19][49] , 
    \couts[19][48] , \couts[19][47] , \couts[19][46] , \couts[19][45] , \couts[19][44] , 
    \couts[19][43] , \couts[19][42] , \couts[19][41] , \couts[19][40] , \couts[19][39] , 
    \couts[19][38] , \couts[19][37] , \couts[19][36] , \couts[19][35] , \couts[19][34] , 
    \couts[19][33] , \couts[19][32] , \couts[19][31] , \couts[19][30] , \couts[19][29] , 
    \couts[19][28] , \couts[19][27] , \couts[19][26] , \couts[19][25] , \couts[19][24] , 
    \couts[19][23] , \couts[19][22] , \couts[19][21] , \couts[19][20] , \couts[19][19] , 
    \couts[19][18] , \couts[19][17] , uc_3211, uc_3212, uc_3213, uc_3214, uc_3215, 
    uc_3216, uc_3217, uc_3218, uc_3219, uc_3220, uc_3221, uc_3222, uc_3223, uc_3224, 
    uc_3225, uc_3226, uc_3227}));
CSA__4_8 CSA19 (.u ({\sums[19][63] , uc_3116, uc_3117, uc_3118, uc_3119, uc_3120, 
    uc_3121, uc_3122, uc_3123, uc_3124, \sums[19][53] , \sums[19][52] , \sums[19][51] , 
    \sums[19][50] , \sums[19][49] , \sums[19][48] , \sums[19][47] , \sums[19][46] , 
    \sums[19][45] , \sums[19][44] , \sums[19][43] , \sums[19][42] , \sums[19][41] , 
    \sums[19][40] , \sums[19][39] , \sums[19][38] , \sums[19][37] , \sums[19][36] , 
    \sums[19][35] , \sums[19][34] , \sums[19][33] , \sums[19][32] , \sums[19][31] , 
    \sums[19][30] , \sums[19][29] , \sums[19][28] , \sums[19][27] , \sums[19][26] , 
    \sums[19][25] , \sums[19][24] , \sums[19][23] , \sums[19][22] , \sums[19][21] , 
    \sums[19][20] , \sums[19][19] , \sums[19][18] , \sums[19][17] , \sums[19][16] , 
    uc_3125, uc_3126, uc_3127, uc_3128, uc_3129, uc_3130, uc_3131, uc_3132, uc_3133, 
    uc_3134, uc_3135, uc_3136, uc_3137, uc_3138, uc_3139, uc_3140}), .v ({\couts[19][63] , 
    uc_3141, uc_3142, uc_3143, uc_3144, uc_3145, uc_3146, uc_3147, uc_3148, \couts[19][54] , 
    \couts[19][53] , \couts[19][52] , \couts[19][51] , \couts[19][50] , \couts[19][49] , 
    \couts[19][48] , \couts[19][47] , \couts[19][46] , \couts[19][45] , \couts[19][44] , 
    \couts[19][43] , \couts[19][42] , \couts[19][41] , \couts[19][40] , \couts[19][39] , 
    \couts[19][38] , \couts[19][37] , \couts[19][36] , \couts[19][35] , \couts[19][34] , 
    \couts[19][33] , \couts[19][32] , \couts[19][31] , \couts[19][30] , \couts[19][29] , 
    \couts[19][28] , \couts[19][27] , \couts[19][26] , \couts[19][25] , \couts[19][24] , 
    \couts[19][23] , \couts[19][22] , \couts[19][21] , \couts[19][20] , \couts[19][19] , 
    \couts[19][18] , \couts[19][17] , uc_3149, uc_3150, uc_3151, uc_3152, uc_3153, 
    uc_3154, uc_3155, uc_3156, uc_3157, uc_3158, uc_3159, uc_3160, uc_3161, uc_3162, 
    uc_3163, uc_3164, uc_3165}), .x ({\sums[13][63] , uc_3030, uc_3031, uc_3032, 
    uc_3033, uc_3034, uc_3035, uc_3036, uc_3037, uc_3038, uc_3039, uc_3040, uc_3041, 
    uc_3042, uc_3043, \sums[13][48] , \sums[13][47] , \sums[13][46] , \sums[13][45] , 
    \sums[13][44] , \sums[13][43] , \sums[13][42] , \sums[13][41] , \sums[13][40] , 
    \sums[13][39] , \sums[13][38] , \sums[13][37] , \sums[13][36] , \sums[13][35] , 
    \sums[13][34] , \sums[13][33] , \sums[13][32] , \sums[13][31] , \sums[13][30] , 
    \sums[13][29] , \sums[13][28] , \sums[13][27] , \sums[13][26] , \sums[13][25] , 
    \sums[13][24] , \sums[13][23] , \sums[13][22] , \sums[13][21] , \sums[13][20] , 
    \sums[13][19] , \sums[13][18] , \sums[13][17] , \sums[13][16] , uc_3044, uc_3045, 
    uc_3046, uc_3047, uc_3048, uc_3049, uc_3050, uc_3051, uc_3052, uc_3053, uc_3054, 
    uc_3055, uc_3056, uc_3057, uc_3058, uc_3059}), .y ({\couts[13][63] , uc_3060, 
    uc_3061, uc_3062, uc_3063, uc_3064, uc_3065, uc_3066, uc_3067, uc_3068, uc_3069, 
    uc_3070, uc_3071, uc_3072, \couts[13][49] , \couts[13][48] , \couts[13][47] , 
    \couts[13][46] , \couts[13][45] , \couts[13][44] , \couts[13][43] , \couts[13][42] , 
    \couts[13][41] , \couts[13][40] , \couts[13][39] , \couts[13][38] , \couts[13][37] , 
    \couts[13][36] , \couts[13][35] , \couts[13][34] , \couts[13][33] , \couts[13][32] , 
    \couts[13][31] , \couts[13][30] , \couts[13][29] , \couts[13][28] , \couts[13][27] , 
    \couts[13][26] , \couts[13][25] , \couts[13][24] , \couts[13][23] , \couts[13][22] , 
    \couts[13][21] , \couts[13][20] , \couts[13][19] , \couts[13][18] , \couts[13][17] , 
    \couts[13][16] , uc_3073, uc_3074, uc_3075, uc_3076, uc_3077, uc_3078, uc_3079, 
    uc_3080, uc_3081, uc_3082, uc_3083, uc_3084, uc_3085, uc_3086, uc_3087, uc_3088})
    , .z ({\sums[14][63] , uc_3089, uc_3090, uc_3091, uc_3092, uc_3093, uc_3094, 
    uc_3095, uc_3096, uc_3097, \sums[14][53] , \sums[14][52] , \sums[14][51] , \sums[14][50] , 
    \sums[14][49] , \sums[14][48] , \sums[14][47] , \sums[14][46] , \sums[14][45] , 
    \sums[14][44] , \sums[14][43] , \sums[14][42] , \sums[14][41] , \sums[14][40] , 
    \sums[14][39] , \sums[14][38] , \sums[14][37] , \sums[14][36] , \sums[14][35] , 
    \sums[14][34] , \sums[14][33] , \sums[14][32] , \sums[14][31] , \sums[14][30] , 
    \sums[14][29] , \sums[14][28] , \sums[14][27] , \sums[14][26] , \sums[14][25] , 
    \sums[14][24] , \sums[14][23] , \sums[14][22] , \sums[14][21] , \sums[14][20] , 
    \sums[6][19] , \pp[18][18] , uc_3098, uc_3099, uc_3100, uc_3101, uc_3102, uc_3103, 
    uc_3104, uc_3105, uc_3106, uc_3107, uc_3108, uc_3109, uc_3110, uc_3111, uc_3112, 
    uc_3113, uc_3114, uc_3115}));
CSA__4_5 CSA14 (.u ({\sums[14][63] , uc_2972, uc_2973, uc_2974, uc_2975, uc_2976, 
    uc_2977, uc_2978, uc_2979, uc_2980, \sums[14][53] , \sums[14][52] , \sums[14][51] , 
    \sums[14][50] , \sums[14][49] , \sums[14][48] , \sums[14][47] , \sums[14][46] , 
    \sums[14][45] , \sums[14][44] , \sums[14][43] , \sums[14][42] , \sums[14][41] , 
    \sums[14][40] , \sums[14][39] , \sums[14][38] , \sums[14][37] , \sums[14][36] , 
    \sums[14][35] , \sums[14][34] , \sums[14][33] , \sums[14][32] , \sums[14][31] , 
    \sums[14][30] , \sums[14][29] , \sums[14][28] , \sums[14][27] , \sums[14][26] , 
    \sums[14][25] , \sums[14][24] , \sums[14][23] , \sums[14][22] , \sums[14][21] , 
    \sums[14][20] , uc_2981, uc_2982, uc_2983, uc_2984, uc_2985, uc_2986, uc_2987, 
    uc_2988, uc_2989, uc_2990, uc_2991, uc_2992, uc_2993, uc_2994, uc_2995, uc_2996, 
    uc_2997, uc_2998, uc_2999, uc_3000}), .v ({\couts[14][63] , uc_3001, uc_3002, 
    uc_3003, uc_3004, uc_3005, uc_3006, uc_3007, uc_3008, \couts[14][54] , \couts[14][53] , 
    \couts[14][52] , \couts[14][51] , \couts[14][50] , \couts[14][49] , \couts[14][48] , 
    \couts[14][47] , \couts[14][46] , \couts[14][45] , \couts[14][44] , \couts[14][43] , 
    \couts[14][42] , \couts[14][41] , \couts[14][40] , \couts[14][39] , \couts[14][38] , 
    \couts[14][37] , \couts[14][36] , \couts[14][35] , \couts[14][34] , \couts[14][33] , 
    \couts[14][32] , \couts[14][31] , \couts[14][30] , \couts[14][29] , \couts[14][28] , 
    \couts[14][27] , \couts[14][26] , \couts[14][25] , \couts[14][24] , \couts[14][23] , 
    \sums[20][22] , \sums[20][21] , uc_3009, uc_3010, uc_3011, uc_3012, uc_3013, 
    uc_3014, uc_3015, uc_3016, uc_3017, uc_3018, uc_3019, uc_3020, uc_3021, uc_3022, 
    uc_3023, uc_3024, uc_3025, uc_3026, uc_3027, uc_3028, uc_3029}), .x ({\sums[6][63] , 
    uc_2879, uc_2880, uc_2881, uc_2882, uc_2883, uc_2884, uc_2885, uc_2886, uc_2887, 
    uc_2888, uc_2889, uc_2890, \sums[6][50] , \sums[6][49] , \sums[6][48] , \sums[6][47] , 
    \sums[6][46] , \sums[6][45] , \sums[6][44] , \sums[6][43] , \sums[6][42] , \sums[6][41] , 
    \sums[6][40] , \sums[6][39] , \sums[6][38] , \sums[6][37] , \sums[6][36] , \sums[6][35] , 
    \sums[6][34] , \sums[6][33] , \sums[6][32] , \sums[6][31] , \sums[6][30] , \sums[6][29] , 
    \sums[6][28] , \sums[6][27] , \sums[6][26] , \sums[6][25] , \sums[6][24] , \sums[6][23] , 
    \sums[6][22] , \sums[6][21] , \sums[6][20] , uc_2891, uc_2892, uc_2893, uc_2894, 
    uc_2895, uc_2896, uc_2897, uc_2898, uc_2899, uc_2900, uc_2901, uc_2902, uc_2903, 
    uc_2904, uc_2905, uc_2906, uc_2907, uc_2908, uc_2909, uc_2910}), .y ({\couts[6][63] , 
    uc_2911, uc_2912, uc_2913, uc_2914, uc_2915, uc_2916, uc_2917, uc_2918, uc_2919, 
    uc_2920, uc_2921, \couts[6][51] , \couts[6][50] , \couts[6][49] , \couts[6][48] , 
    \couts[6][47] , \couts[6][46] , \couts[6][45] , \couts[6][44] , \couts[6][43] , 
    \couts[6][42] , \couts[6][41] , \couts[6][40] , \couts[6][39] , \couts[6][38] , 
    \couts[6][37] , \couts[6][36] , \couts[6][35] , \couts[6][34] , \couts[6][33] , 
    \couts[6][32] , \couts[6][31] , \couts[6][30] , \couts[6][29] , \couts[6][28] , 
    \couts[6][27] , \couts[6][26] , \couts[6][25] , \couts[6][24] , \couts[6][23] , 
    \couts[6][22] , \couts[6][21] , \couts[6][20] , uc_2922, uc_2923, uc_2924, uc_2925, 
    uc_2926, uc_2927, uc_2928, uc_2929, uc_2930, uc_2931, uc_2932, uc_2933, uc_2934, 
    uc_2935, uc_2936, uc_2937, uc_2938, uc_2939, uc_2940, uc_2941}), .z ({\sums[7][63] , 
    uc_2942, uc_2943, uc_2944, uc_2945, uc_2946, uc_2947, uc_2948, uc_2949, uc_2950, 
    \sums[7][53] , \sums[7][52] , \sums[7][51] , \sums[7][50] , \sums[7][49] , \sums[7][48] , 
    \sums[7][47] , \sums[7][46] , \sums[7][45] , \sums[7][44] , \sums[7][43] , \sums[7][42] , 
    \sums[7][41] , \sums[7][40] , \sums[7][39] , \sums[7][38] , \sums[7][37] , \sums[7][36] , 
    \sums[7][35] , \sums[7][34] , \sums[7][33] , \sums[7][32] , \sums[7][31] , \sums[7][30] , 
    \sums[7][29] , \sums[7][28] , \sums[7][27] , \sums[7][26] , \sums[7][25] , \sums[7][24] , 
    \sums[7][23] , \sums[7][22] , \pp[21][21] , uc_2951, uc_2952, uc_2953, uc_2954, 
    uc_2955, uc_2956, uc_2957, uc_2958, uc_2959, uc_2960, uc_2961, uc_2962, uc_2963, 
    uc_2964, uc_2965, uc_2966, uc_2967, uc_2968, uc_2969, uc_2970, uc_2971}));
CSA__4_2 CSA7 (.u ({\sums[7][63] , uc_2817, uc_2818, uc_2819, uc_2820, uc_2821, uc_2822, 
    uc_2823, uc_2824, uc_2825, \sums[7][53] , \sums[7][52] , \sums[7][51] , \sums[7][50] , 
    \sums[7][49] , \sums[7][48] , \sums[7][47] , \sums[7][46] , \sums[7][45] , \sums[7][44] , 
    \sums[7][43] , \sums[7][42] , \sums[7][41] , \sums[7][40] , \sums[7][39] , \sums[7][38] , 
    \sums[7][37] , \sums[7][36] , \sums[7][35] , \sums[7][34] , \sums[7][33] , \sums[7][32] , 
    \sums[7][31] , \sums[7][30] , \sums[7][29] , \sums[7][28] , \sums[7][27] , \sums[7][26] , 
    \sums[7][25] , \sums[7][24] , \sums[7][23] , \sums[7][22] , uc_2826, uc_2827, 
    uc_2828, uc_2829, uc_2830, uc_2831, uc_2832, uc_2833, uc_2834, uc_2835, uc_2836, 
    uc_2837, uc_2838, uc_2839, uc_2840, uc_2841, uc_2842, uc_2843, uc_2844, uc_2845, 
    uc_2846, uc_2847}), .v ({\couts[7][63] , uc_2848, uc_2849, uc_2850, uc_2851, 
    uc_2852, uc_2853, uc_2854, uc_2855, \couts[7][54] , \couts[7][53] , \couts[7][52] , 
    \couts[7][51] , \couts[7][50] , \couts[7][49] , \couts[7][48] , \couts[7][47] , 
    \couts[7][46] , \couts[7][45] , \couts[7][44] , \couts[7][43] , \couts[7][42] , 
    \couts[7][41] , \couts[7][40] , \couts[7][39] , \couts[7][38] , \couts[7][37] , 
    \couts[7][36] , \couts[7][35] , \couts[7][34] , \couts[7][33] , \couts[7][32] , 
    \couts[7][31] , \couts[7][30] , \couts[7][29] , \couts[7][28] , \couts[7][27] , 
    \couts[7][26] , \couts[7][25] , \couts[7][24] , \couts[7][23] , uc_2856, uc_2857, 
    uc_2858, uc_2859, uc_2860, uc_2861, uc_2862, uc_2863, uc_2864, uc_2865, uc_2866, 
    uc_2867, uc_2868, uc_2869, uc_2870, uc_2871, uc_2872, uc_2873, uc_2874, uc_2875, 
    uc_2876, uc_2877, uc_2878}), .x ({\pp[21][63] , uc_2720, uc_2721, uc_2722, uc_2723, 
    uc_2724, uc_2725, uc_2726, uc_2727, uc_2728, uc_2729, uc_2730, \pp[21][51] , 
    \pp[21][50] , \pp[21][49] , \pp[21][48] , \pp[21][47] , \pp[21][46] , \pp[21][45] , 
    \pp[21][44] , \pp[21][43] , \pp[21][42] , \pp[21][41] , \pp[21][40] , \pp[21][39] , 
    \pp[21][38] , \pp[21][37] , \pp[21][36] , \pp[21][35] , \pp[21][34] , \pp[21][33] , 
    \pp[21][32] , \pp[21][31] , \pp[21][30] , \pp[21][29] , \pp[21][28] , \pp[21][27] , 
    \pp[21][26] , \pp[21][25] , \pp[21][24] , \pp[21][23] , \pp[21][22] , uc_2731, 
    uc_2732, uc_2733, uc_2734, uc_2735, uc_2736, uc_2737, uc_2738, uc_2739, uc_2740, 
    uc_2741, uc_2742, uc_2743, uc_2744, uc_2745, uc_2746, uc_2747, uc_2748, uc_2749, 
    uc_2750, uc_2751, uc_2752}), .y ({\pp[22][63] , uc_2753, uc_2754, uc_2755, uc_2756, 
    uc_2757, uc_2758, uc_2759, uc_2760, uc_2761, uc_2762, \pp[22][52] , \pp[22][51] , 
    \pp[22][50] , \pp[22][49] , \pp[22][48] , \pp[22][47] , \pp[22][46] , \pp[22][45] , 
    \pp[22][44] , \pp[22][43] , \pp[22][42] , \pp[22][41] , \pp[22][40] , \pp[22][39] , 
    \pp[22][38] , \pp[22][37] , \pp[22][36] , \pp[22][35] , \pp[22][34] , \pp[22][33] , 
    \pp[22][32] , \pp[22][31] , \pp[22][30] , \pp[22][29] , \pp[22][28] , \pp[22][27] , 
    \pp[22][26] , \pp[22][25] , \pp[22][24] , \pp[22][23] , \pp[22][22] , uc_2763, 
    uc_2764, uc_2765, uc_2766, uc_2767, uc_2768, uc_2769, uc_2770, uc_2771, uc_2772, 
    uc_2773, uc_2774, uc_2775, uc_2776, uc_2777, uc_2778, uc_2779, uc_2780, uc_2781, 
    uc_2782, uc_2783, uc_2784}), .z ({\pp[23][63] , uc_2785, uc_2786, uc_2787, uc_2788, 
    uc_2789, uc_2790, uc_2791, uc_2792, uc_2793, \pp[23][53] , \pp[23][52] , \pp[23][51] , 
    \pp[23][50] , \pp[23][49] , \pp[23][48] , \pp[23][47] , \pp[23][46] , \pp[23][45] , 
    \pp[23][44] , \pp[23][43] , \pp[23][42] , \pp[23][41] , \pp[23][40] , \pp[23][39] , 
    \pp[23][38] , \pp[23][37] , \pp[23][36] , \pp[23][35] , \pp[23][34] , \pp[23][33] , 
    \pp[23][32] , \pp[23][31] , \pp[23][30] , \pp[23][29] , \pp[23][28] , \pp[23][27] , 
    \pp[23][26] , \pp[23][25] , \pp[23][24] , \pp[23][23] , uc_2794, uc_2795, uc_2796, 
    uc_2797, uc_2798, uc_2799, uc_2800, uc_2801, uc_2802, uc_2803, uc_2804, uc_2805, 
    uc_2806, uc_2807, uc_2808, uc_2809, uc_2810, uc_2811, uc_2812, uc_2813, uc_2814, 
    uc_2815, uc_2816}));
CSA__0_75 CSA25 (.u ({\sums[25][63] , \sums[25][62] , \sums[25][61] , \sums[25][60] , 
    \sums[25][59] , \sums[25][58] , \sums[25][57] , \sums[25][56] , \sums[25][55] , 
    \sums[25][54] , \sums[25][53] , \sums[25][52] , \sums[25][51] , \sums[25][50] , 
    \sums[25][49] , \sums[25][48] , \sums[25][47] , \sums[25][46] , \sums[25][45] , 
    \sums[25][44] , \sums[25][43] , \sums[25][42] , \sums[25][41] , \sums[25][40] , 
    \sums[25][39] , \sums[25][38] , \sums[25][37] , \sums[25][36] , \sums[25][35] , 
    \sums[25][34] , \sums[25][33] , \sums[25][32] , \sums[25][31] , \sums[25][30] , 
    \sums[25][29] , \sums[25][28] , \sums[25][27] , \sums[25][26] , \sums[25][25] , 
    \sums[25][24] , \sums[25][23] , \sums[25][22] , \sums[25][21] , \sums[25][20] , 
    \sums[25][19] , \sums[25][18] , \sums[25][17] , \sums[25][16] , \sums[25][15] , 
    \sums[25][14] , \sums[25][13] , \sums[25][12] , \sums[25][11] , \sums[25][10] , 
    \sums[25][9] , \sums[25][8] , \sums[25][7] , \sums[25][6] , out[5], uc_2709, 
    uc_2710, uc_2711, uc_2712, uc_2713}), .v ({\couts[25][63] , \couts[25][62] , 
    \couts[25][61] , \couts[25][60] , \couts[25][59] , \couts[25][58] , \couts[25][57] , 
    \couts[25][56] , \couts[25][55] , \couts[25][54] , \couts[25][53] , \couts[25][52] , 
    \couts[25][51] , \couts[25][50] , \couts[25][49] , \couts[25][48] , \couts[25][47] , 
    \couts[25][46] , \couts[25][45] , \couts[25][44] , \couts[25][43] , \couts[25][42] , 
    \couts[25][41] , \couts[25][40] , \couts[25][39] , \couts[25][38] , \couts[25][37] , 
    \couts[25][36] , \couts[25][35] , \couts[25][34] , \couts[25][33] , \couts[25][32] , 
    \couts[25][31] , \couts[25][30] , \couts[25][29] , \couts[25][28] , \couts[25][27] , 
    \couts[25][26] , \couts[25][25] , \couts[25][24] , \couts[25][23] , \couts[25][22] , 
    \couts[25][21] , \couts[25][20] , \couts[25][19] , \couts[25][18] , \couts[25][17] , 
    \couts[25][16] , \couts[25][15] , \couts[25][14] , \couts[25][13] , \couts[25][12] , 
    \couts[25][11] , \couts[25][10] , \couts[25][9] , \couts[25][8] , \couts[25][7] , 
    \couts[25][6] , uc_2714, uc_2715, uc_2716, uc_2717, uc_2718, uc_2719}), .x ({
    \sums[22][63] , \sums[22][62] , \sums[22][61] , \sums[22][60] , \sums[22][59] , 
    \sums[22][58] , \sums[22][57] , \sums[22][56] , \sums[22][55] , \sums[22][54] , 
    \sums[22][53] , \sums[22][52] , \sums[22][51] , \sums[22][50] , \sums[22][49] , 
    \sums[22][48] , \sums[22][47] , \sums[22][46] , \sums[22][45] , \sums[22][44] , 
    \sums[22][43] , \sums[22][42] , \sums[22][41] , \sums[22][40] , \sums[22][39] , 
    \sums[22][38] , \sums[22][37] , \sums[22][36] , \sums[22][35] , \sums[22][34] , 
    \sums[22][33] , \sums[22][32] , \sums[22][31] , \sums[22][30] , \sums[22][29] , 
    \sums[22][28] , \sums[22][27] , \sums[22][26] , \sums[22][25] , \sums[22][24] , 
    \sums[22][23] , \sums[22][22] , \sums[22][21] , \sums[22][20] , \sums[22][19] , 
    \sums[22][18] , \sums[22][17] , \sums[22][16] , \sums[22][15] , \sums[22][14] , 
    \sums[22][13] , \sums[22][12] , \sums[22][11] , \sums[22][10] , \sums[22][9] , 
    \sums[22][8] , \sums[22][7] , \sums[22][6] , \sums[22][5] , uc_2689, uc_2690, 
    uc_2691, uc_2692, uc_2693}), .y ({\couts[22][63] , \couts[22][62] , \couts[22][61] , 
    \couts[22][60] , \couts[22][59] , \couts[22][58] , \couts[22][57] , \couts[22][56] , 
    \couts[22][55] , \couts[22][54] , \couts[22][53] , \couts[22][52] , \couts[22][51] , 
    \couts[22][50] , \couts[22][49] , \couts[22][48] , \couts[22][47] , \couts[22][46] , 
    \couts[22][45] , \couts[22][44] , \couts[22][43] , \couts[22][42] , \couts[22][41] , 
    \couts[22][40] , \couts[22][39] , \couts[22][38] , \couts[22][37] , \couts[22][36] , 
    \couts[22][35] , \couts[22][34] , \couts[22][33] , \couts[22][32] , \couts[22][31] , 
    \couts[22][30] , \couts[22][29] , \couts[22][28] , \couts[22][27] , \couts[22][26] , 
    \couts[22][25] , \couts[22][24] , \couts[22][23] , \couts[22][22] , \couts[22][21] , 
    \couts[22][20] , \couts[22][19] , \couts[22][18] , \couts[22][17] , \couts[22][16] , 
    \couts[22][15] , \couts[22][14] , \couts[22][13] , \couts[22][12] , \couts[22][11] , 
    \couts[22][10] , \couts[22][9] , \couts[22][8] , \couts[22][7] , \couts[22][6] , 
    \couts[22][5] , uc_2694, uc_2695, uc_2696, uc_2697, uc_2698}), .z ({\sums[23][63] , 
    \sums[23][62] , \sums[23][61] , \sums[23][60] , \sums[23][59] , \sums[23][58] , 
    \sums[23][57] , \sums[23][56] , \sums[23][55] , \sums[23][54] , \sums[23][53] , 
    \sums[23][52] , \sums[23][51] , \sums[23][50] , \sums[23][49] , \sums[23][48] , 
    \sums[23][47] , \sums[23][46] , \sums[23][45] , \sums[23][44] , \sums[23][43] , 
    \sums[23][42] , \sums[23][41] , \sums[23][40] , \sums[23][39] , \sums[23][38] , 
    \sums[23][37] , \sums[23][36] , \sums[23][35] , \sums[23][34] , \sums[23][33] , 
    \sums[23][32] , \sums[23][31] , \sums[23][30] , \sums[23][29] , \sums[23][28] , 
    \sums[23][27] , \sums[23][26] , \sums[23][25] , \sums[23][24] , \sums[23][23] , 
    \sums[23][22] , \sums[23][21] , \sums[23][20] , \sums[23][19] , \sums[23][18] , 
    \sums[23][17] , \sums[23][16] , \sums[23][15] , \sums[23][14] , \couts[18][13] , 
    \couts[18][12] , \couts[18][11] , \couts[18][10] , uc_2699, uc_2700, uc_2701, 
    uc_2702, uc_2703, uc_2704, uc_2705, uc_2706, uc_2707, uc_2708}));
CSA__3_14 CSA0 (.u ({uc_2627, uc_2628, \sums[0][61] , uc_2629, uc_2630, uc_2631, 
    uc_2632, uc_2633, uc_2634, uc_2635, uc_2636, uc_2637, uc_2638, uc_2639, uc_2640, 
    uc_2641, uc_2642, uc_2643, uc_2644, uc_2645, uc_2646, uc_2647, uc_2648, uc_2649, 
    uc_2650, uc_2651, uc_2652, uc_2653, uc_2654, uc_2655, uc_2656, \sums[0][32] , 
    \sums[0][31] , \sums[0][30] , \sums[0][29] , \sums[0][28] , \sums[0][27] , \sums[0][26] , 
    \sums[0][25] , \sums[0][24] , \sums[0][23] , \sums[0][22] , \sums[0][21] , \sums[0][20] , 
    \sums[0][19] , \sums[0][18] , \sums[0][17] , \sums[0][16] , \sums[0][15] , \sums[0][14] , 
    \sums[0][13] , \sums[0][12] , \sums[0][11] , \sums[0][10] , \sums[0][9] , \sums[0][8] , 
    \sums[0][7] , \sums[0][6] , \sums[0][5] , \sums[0][4] , \sums[0][3] , \sums[0][2] , 
    out[1], uc_2657}), .v ({uc_2658, uc_2659, \couts[0][61] , uc_2660, uc_2661, uc_2662, 
    uc_2663, uc_2664, uc_2665, uc_2666, uc_2667, uc_2668, uc_2669, uc_2670, uc_2671, 
    uc_2672, uc_2673, uc_2674, uc_2675, uc_2676, uc_2677, uc_2678, uc_2679, uc_2680, 
    uc_2681, uc_2682, uc_2683, uc_2684, uc_2685, uc_2686, \couts[0][33] , \couts[0][32] , 
    \couts[0][31] , \couts[0][30] , \couts[0][29] , \couts[0][28] , \couts[0][27] , 
    \couts[0][26] , \couts[0][25] , \couts[0][24] , \couts[0][23] , \couts[0][22] , 
    \couts[0][21] , \couts[0][20] , \couts[0][19] , \couts[0][18] , \couts[0][17] , 
    \couts[0][16] , \couts[0][15] , \couts[0][14] , \couts[0][13] , \couts[0][12] , 
    \couts[0][11] , \couts[0][10] , \couts[0][9] , \couts[0][8] , \couts[0][7] , 
    \couts[0][6] , \couts[0][5] , \couts[0][4] , \couts[0][3] , \couts[0][2] , uc_2687, 
    uc_2688}), .x ({uc_2530, uc_2531, \pp[0][63] , uc_2532, uc_2533, uc_2534, uc_2535, 
    uc_2536, uc_2537, uc_2538, uc_2539, uc_2540, uc_2541, uc_2542, uc_2543, uc_2544, 
    uc_2545, uc_2546, uc_2547, uc_2548, uc_2549, uc_2550, uc_2551, uc_2552, uc_2553, 
    uc_2554, uc_2555, uc_2556, uc_2557, uc_2558, uc_2559, uc_2560, uc_2561, \pp[0][30] , 
    \pp[0][29] , \pp[0][28] , \pp[0][27] , \pp[0][26] , \pp[0][25] , \pp[0][24] , 
    \pp[0][23] , \pp[0][22] , \pp[0][21] , \pp[0][20] , \pp[0][19] , \pp[0][18] , 
    \pp[0][17] , \pp[0][16] , \pp[0][15] , \pp[0][14] , \pp[0][13] , \pp[0][12] , 
    \pp[0][11] , \pp[0][10] , \pp[0][9] , \pp[0][8] , \pp[0][7] , \pp[0][6] , \pp[0][5] , 
    \pp[0][4] , \pp[0][3] , \pp[0][2] , \pp[0][1] , uc_2562}), .y ({uc_2563, uc_2564, 
    \pp[1][63] , uc_2565, uc_2566, uc_2567, uc_2568, uc_2569, uc_2570, uc_2571, uc_2572, 
    uc_2573, uc_2574, uc_2575, uc_2576, uc_2577, uc_2578, uc_2579, uc_2580, uc_2581, 
    uc_2582, uc_2583, uc_2584, uc_2585, uc_2586, uc_2587, uc_2588, uc_2589, uc_2590, 
    uc_2591, uc_2592, uc_2593, \pp[1][31] , \pp[1][30] , \pp[1][29] , \pp[1][28] , 
    \pp[1][27] , \pp[1][26] , \pp[1][25] , \pp[1][24] , \pp[1][23] , \pp[1][22] , 
    \pp[1][21] , \pp[1][20] , \pp[1][19] , \pp[1][18] , \pp[1][17] , \pp[1][16] , 
    \pp[1][15] , \pp[1][14] , \pp[1][13] , \pp[1][12] , \pp[1][11] , \pp[1][10] , 
    \pp[1][9] , \pp[1][8] , \pp[1][7] , \pp[1][6] , \pp[1][5] , \pp[1][4] , \pp[1][3] , 
    \pp[1][2] , \pp[1][1] , uc_2594}), .z ({uc_2595, uc_2596, \pp[2][63] , uc_2597, 
    uc_2598, uc_2599, uc_2600, uc_2601, uc_2602, uc_2603, uc_2604, uc_2605, uc_2606, 
    uc_2607, uc_2608, uc_2609, uc_2610, uc_2611, uc_2612, uc_2613, uc_2614, uc_2615, 
    uc_2616, uc_2617, uc_2618, uc_2619, uc_2620, uc_2621, uc_2622, uc_2623, uc_2624, 
    \pp[2][32] , \pp[2][31] , \pp[2][30] , \pp[2][29] , \pp[2][28] , \pp[2][27] , 
    \pp[2][26] , \pp[2][25] , \pp[2][24] , \pp[2][23] , \pp[2][22] , \pp[2][21] , 
    \pp[2][20] , \pp[2][19] , \pp[2][18] , \pp[2][17] , \pp[2][16] , \pp[2][15] , 
    \pp[2][14] , \pp[2][13] , \pp[2][12] , \pp[2][11] , \pp[2][10] , \pp[2][9] , 
    \pp[2][8] , \pp[2][7] , \pp[2][6] , \pp[2][5] , \pp[2][4] , \pp[2][3] , \pp[2][2] , 
    uc_2625, uc_2626}));
CSA__3_11 CSA1 (.u ({uc_2468, uc_2469, \sums[1][61] , uc_2470, uc_2471, uc_2472, 
    uc_2473, uc_2474, uc_2475, uc_2476, uc_2477, uc_2478, uc_2479, uc_2480, uc_2481, 
    uc_2482, uc_2483, uc_2484, uc_2485, uc_2486, uc_2487, uc_2488, uc_2489, uc_2490, 
    uc_2491, uc_2492, uc_2493, uc_2494, \sums[1][35] , \sums[1][34] , \sums[1][33] , 
    \sums[1][32] , \sums[1][31] , \sums[1][30] , \sums[1][29] , \sums[1][28] , \sums[1][27] , 
    \sums[1][26] , \sums[1][25] , \sums[1][24] , \sums[1][23] , \sums[1][22] , \sums[1][21] , 
    \sums[1][20] , \sums[1][19] , \sums[1][18] , \sums[1][17] , \sums[1][16] , \sums[1][15] , 
    \sums[1][14] , \sums[1][13] , \sums[1][12] , \sums[1][11] , \sums[1][10] , \sums[1][9] , 
    \sums[1][8] , \sums[1][7] , \sums[1][6] , \sums[1][5] , \sums[1][4] , uc_2495, 
    uc_2496, uc_2497, uc_2498}), .v ({\couts[1][37] , uc_2499, uc_2500, uc_2501, 
    uc_2502, uc_2503, uc_2504, uc_2505, uc_2506, uc_2507, uc_2508, uc_2509, uc_2510, 
    uc_2511, uc_2512, uc_2513, uc_2514, uc_2515, uc_2516, uc_2517, uc_2518, uc_2519, 
    uc_2520, uc_2521, uc_2522, uc_2523, uc_2524, \couts[1][36] , \couts[1][35] , 
    \couts[1][34] , \couts[1][33] , \couts[1][32] , \couts[1][31] , \couts[1][30] , 
    \couts[1][29] , \couts[1][28] , \couts[1][27] , \couts[1][26] , \couts[1][25] , 
    \couts[1][24] , \couts[1][23] , \couts[1][22] , \couts[1][21] , \couts[1][20] , 
    \couts[1][19] , \couts[1][18] , \couts[1][17] , \couts[1][16] , \couts[1][15] , 
    \couts[1][14] , \couts[1][13] , \couts[1][12] , \couts[1][11] , \couts[1][10] , 
    \couts[1][9] , \couts[1][8] , \couts[1][7] , \couts[1][6] , n_2_0, uc_2525, uc_2526, 
    uc_2527, uc_2528, uc_2529}), .x ({uc_2371, \pp[3][63] , uc_2372, uc_2373, uc_2374, 
    uc_2375, uc_2376, uc_2377, uc_2378, uc_2379, uc_2380, uc_2381, uc_2382, uc_2383, 
    uc_2384, uc_2385, uc_2386, uc_2387, uc_2388, uc_2389, uc_2390, uc_2391, uc_2392, 
    uc_2393, uc_2394, uc_2395, uc_2396, uc_2397, uc_2398, uc_2399, \pp[3][33] , \pp[3][32] , 
    \pp[3][31] , \pp[3][30] , \pp[3][29] , \pp[3][28] , \pp[3][27] , \pp[3][26] , 
    \pp[3][25] , \pp[3][24] , \pp[3][23] , \pp[3][22] , \pp[3][21] , \pp[3][20] , 
    \pp[3][19] , \pp[3][18] , \pp[3][17] , \pp[3][16] , \pp[3][15] , \pp[3][14] , 
    \pp[3][13] , \pp[3][12] , \pp[3][11] , \pp[3][10] , \pp[3][9] , \pp[3][8] , \pp[3][7] , 
    \pp[3][6] , \pp[3][5] , \pp[3][4] , uc_2400, uc_2401, uc_2402, uc_2403}), .y ({
    uc_2404, \pp[4][63] , uc_2405, uc_2406, uc_2407, uc_2408, uc_2409, uc_2410, uc_2411, 
    uc_2412, uc_2413, uc_2414, uc_2415, uc_2416, uc_2417, uc_2418, uc_2419, uc_2420, 
    uc_2421, uc_2422, uc_2423, uc_2424, uc_2425, uc_2426, uc_2427, uc_2428, uc_2429, 
    uc_2430, uc_2431, \pp[4][34] , \pp[4][33] , \pp[4][32] , \pp[4][31] , \pp[4][30] , 
    \pp[4][29] , \pp[4][28] , \pp[4][27] , \pp[4][26] , \pp[4][25] , \pp[4][24] , 
    \pp[4][23] , \pp[4][22] , \pp[4][21] , \pp[4][20] , \pp[4][19] , \pp[4][18] , 
    \pp[4][17] , \pp[4][16] , \pp[4][15] , \pp[4][14] , \pp[4][13] , \pp[4][12] , 
    \pp[4][11] , \pp[4][10] , \pp[4][9] , \pp[4][8] , \pp[4][7] , \pp[4][6] , \pp[4][5] , 
    \pp[4][4] , uc_2432, uc_2433, uc_2434, uc_2435}), .z ({uc_2436, \pp[5][63] , 
    uc_2437, uc_2438, uc_2439, uc_2440, uc_2441, uc_2442, uc_2443, uc_2444, uc_2445, 
    uc_2446, uc_2447, uc_2448, uc_2449, uc_2450, uc_2451, uc_2452, uc_2453, uc_2454, 
    uc_2455, uc_2456, uc_2457, uc_2458, uc_2459, uc_2460, uc_2461, uc_2462, \pp[5][35] , 
    \pp[5][34] , \pp[5][33] , \pp[5][32] , \pp[5][31] , \pp[5][30] , \pp[5][29] , 
    \pp[5][28] , \pp[5][27] , \pp[5][26] , \pp[5][25] , \pp[5][24] , \pp[5][23] , 
    \pp[5][22] , \pp[5][21] , \pp[5][20] , \pp[5][19] , \pp[5][18] , \pp[5][17] , 
    \pp[5][16] , \pp[5][15] , \pp[5][14] , \pp[5][13] , \pp[5][12] , \pp[5][11] , 
    \pp[5][10] , \pp[5][9] , \pp[5][8] , \pp[5][7] , \pp[5][6] , \pp[5][5] , uc_2463, 
    uc_2464, uc_2465, uc_2466, uc_2467}));
CSA__3_8 CSA22 (.u ({\sums[22][63] , \sums[22][62] , \sums[22][61] , \sums[22][60] , 
    \sums[22][59] , \sums[22][58] , \sums[22][57] , \sums[22][56] , \sums[22][55] , 
    \sums[22][54] , \sums[22][53] , \sums[22][52] , \sums[22][51] , \sums[22][50] , 
    \sums[22][49] , \sums[22][48] , \sums[22][47] , \sums[22][46] , \sums[22][45] , 
    \sums[22][44] , \sums[22][43] , \sums[22][42] , \sums[22][41] , \sums[22][40] , 
    \sums[22][39] , \sums[22][38] , \sums[22][37] , \sums[22][36] , \sums[22][35] , 
    \sums[22][34] , \sums[22][33] , \sums[22][32] , \sums[22][31] , \sums[22][30] , 
    \sums[22][29] , \sums[22][28] , \sums[22][27] , \sums[22][26] , \sums[22][25] , 
    \sums[22][24] , \sums[22][23] , \sums[22][22] , \sums[22][21] , \sums[22][20] , 
    \sums[22][19] , \sums[22][18] , \sums[22][17] , \sums[22][16] , \sums[22][15] , 
    \sums[22][14] , \sums[22][13] , \sums[22][12] , \sums[22][11] , \sums[22][10] , 
    \sums[22][9] , \sums[22][8] , \sums[22][7] , \sums[22][6] , \sums[22][5] , out[4], 
    uc_2362, uc_2363, uc_2364, uc_2365}), .v ({\couts[22][63] , \couts[22][62] , 
    \couts[22][61] , \couts[22][60] , \couts[22][59] , \couts[22][58] , \couts[22][57] , 
    \couts[22][56] , \couts[22][55] , \couts[22][54] , \couts[22][53] , \couts[22][52] , 
    \couts[22][51] , \couts[22][50] , \couts[22][49] , \couts[22][48] , \couts[22][47] , 
    \couts[22][46] , \couts[22][45] , \couts[22][44] , \couts[22][43] , \couts[22][42] , 
    \couts[22][41] , \couts[22][40] , \couts[22][39] , \couts[22][38] , \couts[22][37] , 
    \couts[22][36] , \couts[22][35] , \couts[22][34] , \couts[22][33] , \couts[22][32] , 
    \couts[22][31] , \couts[22][30] , \couts[22][29] , \couts[22][28] , \couts[22][27] , 
    \couts[22][26] , \couts[22][25] , \couts[22][24] , \couts[22][23] , \couts[22][22] , 
    \couts[22][21] , \couts[22][20] , \couts[22][19] , \couts[22][18] , \couts[22][17] , 
    \couts[22][16] , \couts[22][15] , \couts[22][14] , \couts[22][13] , \couts[22][12] , 
    \couts[22][11] , \couts[22][10] , \couts[22][9] , \couts[22][8] , \couts[22][7] , 
    \couts[22][6] , \couts[22][5] , uc_2366, uc_2367, uc_2368, uc_2369, uc_2370})
    , .x ({\sums[17][63] , \sums[17][62] , \sums[17][61] , \sums[17][60] , \sums[17][59] , 
    \sums[17][58] , \sums[17][57] , \sums[17][56] , \sums[17][55] , \sums[17][54] , 
    \sums[17][53] , \sums[17][52] , \sums[17][51] , \sums[17][50] , \sums[17][49] , 
    \sums[17][48] , \sums[17][47] , \sums[17][46] , \sums[17][45] , \sums[17][44] , 
    \sums[17][43] , \sums[17][42] , \sums[17][41] , \sums[17][40] , \sums[17][39] , 
    \sums[17][38] , \sums[17][37] , \sums[17][36] , \sums[17][35] , \sums[17][34] , 
    \sums[17][33] , \sums[17][32] , \sums[17][31] , \sums[17][30] , \sums[17][29] , 
    \sums[17][28] , \sums[17][27] , \sums[17][26] , \sums[17][25] , \sums[17][24] , 
    \sums[17][23] , \sums[17][22] , \sums[17][21] , \sums[17][20] , \sums[17][19] , 
    \sums[17][18] , \sums[17][17] , \sums[17][16] , \sums[17][15] , \sums[17][14] , 
    \sums[17][13] , \sums[17][12] , \sums[17][11] , \sums[17][10] , \sums[17][9] , 
    \sums[17][8] , \sums[17][7] , \sums[17][6] , \sums[17][5] , \sums[17][4] , uc_2347, 
    uc_2348, uc_2349, uc_2350}), .y ({\couts[17][63] , \couts[17][62] , \couts[17][61] , 
    \couts[17][60] , \couts[17][59] , \couts[17][58] , \couts[17][57] , \couts[17][56] , 
    \couts[17][55] , \couts[17][54] , \couts[17][53] , \couts[17][52] , \couts[17][51] , 
    \couts[17][50] , \couts[17][49] , \couts[17][48] , \couts[17][47] , \couts[17][46] , 
    \couts[17][45] , \couts[17][44] , \couts[17][43] , \couts[17][42] , \couts[17][41] , 
    \couts[17][40] , \couts[17][39] , \couts[17][38] , \couts[17][37] , \couts[17][36] , 
    \couts[17][35] , \couts[17][34] , \couts[17][33] , \couts[17][32] , \couts[17][31] , 
    \couts[17][30] , \couts[17][29] , \couts[17][28] , \couts[17][27] , \couts[17][26] , 
    \couts[17][25] , \couts[17][24] , \couts[17][23] , \couts[17][22] , \couts[17][21] , 
    \couts[17][20] , \couts[17][19] , \couts[17][18] , \couts[17][17] , \couts[17][16] , 
    \couts[17][15] , \couts[17][14] , \couts[17][13] , \couts[17][12] , \couts[17][11] , 
    \couts[17][10] , \couts[17][9] , \couts[17][8] , \couts[17][7] , \couts[17][6] , 
    \couts[17][5] , \couts[17][4] , uc_2351, uc_2352, uc_2353, uc_2354}), .z ({\sums[18][63] , 
    \sums[18][62] , \sums[18][61] , \sums[18][60] , \sums[18][59] , \sums[18][58] , 
    \sums[18][57] , \sums[18][56] , \sums[18][55] , \sums[18][54] , \sums[18][53] , 
    \sums[18][52] , \sums[18][51] , \sums[18][50] , \sums[18][49] , \sums[18][48] , 
    \sums[18][47] , \sums[18][46] , \sums[18][45] , \sums[18][44] , \sums[18][43] , 
    \sums[18][42] , \sums[18][41] , \sums[18][40] , \sums[18][39] , \sums[18][38] , 
    \sums[18][37] , \sums[18][36] , \sums[18][35] , \sums[18][34] , \sums[18][33] , 
    \sums[18][32] , \sums[18][31] , \sums[18][30] , \sums[18][29] , \sums[18][28] , 
    \sums[18][27] , \sums[18][26] , \sums[18][25] , \sums[18][24] , \sums[18][23] , 
    \sums[18][22] , \sums[18][21] , \sums[18][20] , \sums[18][19] , \sums[18][18] , 
    \sums[18][17] , \sums[18][16] , \sums[18][15] , \sums[18][14] , \sums[18][13] , 
    \sums[18][12] , \sums[18][11] , \sums[18][10] , \sums[18][9] , \sums[18][8] , 
    \sums[18][7] , uc_2355, uc_2356, uc_2357, uc_2358, uc_2359, uc_2360, uc_2361}));
CSA__3_5 CSA10 (.u ({uc_2289, \sums[10][62] , uc_2290, uc_2291, uc_2292, uc_2293, 
    uc_2294, uc_2295, uc_2296, uc_2297, uc_2298, uc_2299, uc_2300, uc_2301, uc_2302, 
    uc_2303, uc_2304, uc_2305, uc_2306, uc_2307, uc_2308, uc_2309, uc_2310, uc_2311, 
    uc_2312, uc_2313, uc_2314, uc_2315, \sums[10][35] , \sums[10][34] , \sums[10][33] , 
    \sums[10][32] , \sums[10][31] , \sums[10][30] , \sums[10][29] , \sums[10][28] , 
    \sums[10][27] , \sums[10][26] , \sums[10][25] , \sums[10][24] , \sums[10][23] , 
    \sums[10][22] , \sums[10][21] , \sums[10][20] , \sums[10][19] , \sums[10][18] , 
    \sums[10][17] , \sums[10][16] , \sums[10][15] , \sums[10][14] , \sums[10][13] , 
    \sums[10][12] , \sums[10][11] , \sums[10][10] , \sums[10][9] , \sums[10][8] , 
    \sums[10][7] , \sums[10][6] , \sums[10][5] , \sums[10][4] , \sums[10][3] , out[2], 
    uc_2316, uc_2317}), .v ({uc_2318, \couts[10][62] , uc_2319, uc_2320, uc_2321, 
    uc_2322, uc_2323, uc_2324, uc_2325, uc_2326, uc_2327, uc_2328, uc_2329, uc_2330, 
    uc_2331, uc_2332, uc_2333, uc_2334, uc_2335, uc_2336, uc_2337, uc_2338, uc_2339, 
    uc_2340, uc_2341, uc_2342, uc_2343, \couts[10][36] , \couts[10][35] , \couts[10][34] , 
    \couts[10][33] , \couts[10][32] , \couts[10][31] , \couts[10][30] , \couts[10][29] , 
    \couts[10][28] , \couts[10][27] , \couts[10][26] , \couts[10][25] , \couts[10][24] , 
    \couts[10][23] , \couts[10][22] , \couts[10][21] , \couts[10][20] , \couts[10][19] , 
    \couts[10][18] , \couts[10][17] , \couts[10][16] , \couts[10][15] , \couts[10][14] , 
    \couts[10][13] , \couts[10][12] , \couts[10][11] , \couts[10][10] , \couts[10][9] , 
    \couts[10][8] , \couts[10][7] , \couts[10][6] , \couts[10][5] , \couts[10][4] , 
    \couts[10][3] , uc_2344, uc_2345, uc_2346}), .x ({uc_2196, uc_2197, \sums[0][61] , 
    uc_2198, uc_2199, uc_2200, uc_2201, uc_2202, uc_2203, uc_2204, uc_2205, uc_2206, 
    uc_2207, uc_2208, uc_2209, uc_2210, uc_2211, uc_2212, uc_2213, uc_2214, uc_2215, 
    uc_2216, uc_2217, uc_2218, uc_2219, uc_2220, uc_2221, uc_2222, uc_2223, uc_2224, 
    uc_2225, \sums[0][32] , \sums[0][31] , \sums[0][30] , \sums[0][29] , \sums[0][28] , 
    \sums[0][27] , \sums[0][26] , \sums[0][25] , \sums[0][24] , \sums[0][23] , \sums[0][22] , 
    \sums[0][21] , \sums[0][20] , \sums[0][19] , \sums[0][18] , \sums[0][17] , \sums[0][16] , 
    \sums[0][15] , \sums[0][14] , \sums[0][13] , \sums[0][12] , \sums[0][11] , \sums[0][10] , 
    \sums[0][9] , \sums[0][8] , \sums[0][7] , \sums[0][6] , \sums[0][5] , \sums[0][4] , 
    \sums[0][3] , \sums[0][2] , uc_2226, uc_2227}), .y ({uc_2228, uc_2229, \couts[0][61] , 
    uc_2230, uc_2231, uc_2232, uc_2233, uc_2234, uc_2235, uc_2236, uc_2237, uc_2238, 
    uc_2239, uc_2240, uc_2241, uc_2242, uc_2243, uc_2244, uc_2245, uc_2246, uc_2247, 
    uc_2248, uc_2249, uc_2250, uc_2251, uc_2252, uc_2253, uc_2254, uc_2255, uc_2256, 
    \couts[0][33] , \couts[0][32] , \couts[0][31] , \couts[0][30] , \couts[0][29] , 
    \couts[0][28] , \couts[0][27] , \couts[0][26] , \couts[0][25] , \couts[0][24] , 
    \couts[0][23] , \couts[0][22] , \couts[0][21] , \couts[0][20] , \couts[0][19] , 
    \couts[0][18] , \couts[0][17] , \couts[0][16] , \couts[0][15] , \couts[0][14] , 
    \couts[0][13] , \couts[0][12] , \couts[0][11] , \couts[0][10] , \couts[0][9] , 
    \couts[0][8] , \couts[0][7] , \couts[0][6] , \couts[0][5] , \couts[0][4] , \couts[0][3] , 
    \couts[0][2] , uc_2257, uc_2258}), .z ({uc_2259, uc_2260, \sums[1][61] , uc_2261, 
    uc_2262, uc_2263, uc_2264, uc_2265, uc_2266, uc_2267, uc_2268, uc_2269, uc_2270, 
    uc_2271, uc_2272, uc_2273, uc_2274, uc_2275, uc_2276, uc_2277, uc_2278, uc_2279, 
    uc_2280, uc_2281, uc_2282, uc_2283, uc_2284, uc_2285, \sums[1][35] , \sums[1][34] , 
    \sums[1][33] , \sums[1][32] , \sums[1][31] , \sums[1][30] , \sums[1][29] , \sums[1][28] , 
    \sums[1][27] , \sums[1][26] , \sums[1][25] , \sums[1][24] , \sums[1][23] , \sums[1][22] , 
    \sums[1][21] , \sums[1][20] , \sums[1][19] , \sums[1][18] , \sums[1][17] , \sums[1][16] , 
    \sums[1][15] , \sums[1][14] , \sums[1][13] , \sums[1][12] , \sums[1][11] , \sums[1][10] , 
    \sums[1][9] , \sums[1][8] , \sums[1][7] , \sums[1][6] , \sums[1][5] , \sums[1][4] , 
    \pp[3][3] , uc_2286, uc_2287, uc_2288}));
CSA__3_2 CSA17 (.u ({\sums[17][63] , \sums[17][62] , \sums[17][61] , \sums[17][60] , 
    \sums[17][59] , \sums[17][58] , \sums[17][57] , \sums[17][56] , \sums[17][55] , 
    \sums[17][54] , \sums[17][53] , \sums[17][52] , \sums[17][51] , \sums[17][50] , 
    \sums[17][49] , \sums[17][48] , \sums[17][47] , \sums[17][46] , \sums[17][45] , 
    \sums[17][44] , \sums[17][43] , \sums[17][42] , \sums[17][41] , \sums[17][40] , 
    \sums[17][39] , \sums[17][38] , \sums[17][37] , \sums[17][36] , \sums[17][35] , 
    \sums[17][34] , \sums[17][33] , \sums[17][32] , \sums[17][31] , \sums[17][30] , 
    \sums[17][29] , \sums[17][28] , \sums[17][27] , \sums[17][26] , \sums[17][25] , 
    \sums[17][24] , \sums[17][23] , \sums[17][22] , \sums[17][21] , \sums[17][20] , 
    \sums[17][19] , \sums[17][18] , \sums[17][17] , \sums[17][16] , \sums[17][15] , 
    \sums[17][14] , \sums[17][13] , \sums[17][12] , \sums[17][11] , \sums[17][10] , 
    \sums[17][9] , \sums[17][8] , \sums[17][7] , \sums[17][6] , \sums[17][5] , \sums[17][4] , 
    out[3], uc_2189, uc_2190, uc_2191}), .v ({\couts[17][63] , \couts[17][62] , \couts[17][61] , 
    \couts[17][60] , \couts[17][59] , \couts[17][58] , \couts[17][57] , \couts[17][56] , 
    \couts[17][55] , \couts[17][54] , \couts[17][53] , \couts[17][52] , \couts[17][51] , 
    \couts[17][50] , \couts[17][49] , \couts[17][48] , \couts[17][47] , \couts[17][46] , 
    \couts[17][45] , \couts[17][44] , \couts[17][43] , \couts[17][42] , \couts[17][41] , 
    \couts[17][40] , \couts[17][39] , \couts[17][38] , \couts[17][37] , \couts[17][36] , 
    \couts[17][35] , \couts[17][34] , \couts[17][33] , \couts[17][32] , \couts[17][31] , 
    \couts[17][30] , \couts[17][29] , \couts[17][28] , \couts[17][27] , \couts[17][26] , 
    \couts[17][25] , \couts[17][24] , \couts[17][23] , \couts[17][22] , \couts[17][21] , 
    \couts[17][20] , \couts[17][19] , \couts[17][18] , \couts[17][17] , \couts[17][16] , 
    \couts[17][15] , \couts[17][14] , \couts[17][13] , \couts[17][12] , \couts[17][11] , 
    \couts[17][10] , \couts[17][9] , \couts[17][8] , \couts[17][7] , \couts[17][6] , 
    \couts[17][5] , \couts[17][4] , uc_2192, uc_2193, uc_2194, uc_2195}), .x ({uc_2125, 
    \sums[10][62] , uc_2126, uc_2127, uc_2128, uc_2129, uc_2130, uc_2131, uc_2132, 
    uc_2133, uc_2134, uc_2135, uc_2136, uc_2137, uc_2138, uc_2139, uc_2140, uc_2141, 
    uc_2142, uc_2143, uc_2144, uc_2145, uc_2146, uc_2147, uc_2148, uc_2149, uc_2150, 
    uc_2151, \sums[10][35] , \sums[10][34] , \sums[10][33] , \sums[10][32] , \sums[10][31] , 
    \sums[10][30] , \sums[10][29] , \sums[10][28] , \sums[10][27] , \sums[10][26] , 
    \sums[10][25] , \sums[10][24] , \sums[10][23] , \sums[10][22] , \sums[10][21] , 
    \sums[10][20] , \sums[10][19] , \sums[10][18] , \sums[10][17] , \sums[10][16] , 
    \sums[10][15] , \sums[10][14] , \sums[10][13] , \sums[10][12] , \sums[10][11] , 
    \sums[10][10] , \sums[10][9] , \sums[10][8] , \sums[10][7] , \sums[10][6] , \sums[10][5] , 
    \sums[10][4] , \sums[10][3] , uc_2152, uc_2153, uc_2154}), .y ({uc_2155, \couts[10][62] , 
    uc_2156, uc_2157, uc_2158, uc_2159, uc_2160, uc_2161, uc_2162, uc_2163, uc_2164, 
    uc_2165, uc_2166, uc_2167, uc_2168, uc_2169, uc_2170, uc_2171, uc_2172, uc_2173, 
    uc_2174, uc_2175, uc_2176, uc_2177, uc_2178, uc_2179, uc_2180, \couts[10][36] , 
    \couts[10][35] , \couts[10][34] , \couts[10][33] , \couts[10][32] , \couts[10][31] , 
    \couts[10][30] , \couts[10][29] , \couts[10][28] , \couts[10][27] , \couts[10][26] , 
    \couts[10][25] , \couts[10][24] , \couts[10][23] , \couts[10][22] , \couts[10][21] , 
    \couts[10][20] , \couts[10][19] , \couts[10][18] , \couts[10][17] , \couts[10][16] , 
    \couts[10][15] , \couts[10][14] , \couts[10][13] , \couts[10][12] , \couts[10][11] , 
    \couts[10][10] , \couts[10][9] , \couts[10][8] , \couts[10][7] , \couts[10][6] , 
    \couts[10][5] , \couts[10][4] , \couts[10][3] , uc_2181, uc_2182, uc_2183}), .z ({
    \sums[11][63] , \sums[11][62] , \sums[11][61] , \sums[11][60] , \sums[11][59] , 
    \sums[11][58] , \sums[11][57] , \sums[11][56] , \sums[11][55] , \sums[11][54] , 
    \sums[11][53] , \sums[11][52] , \sums[11][51] , \sums[11][50] , \sums[11][49] , 
    \sums[11][48] , \sums[11][47] , \sums[11][46] , \sums[11][45] , \sums[11][44] , 
    \sums[11][43] , \sums[11][42] , \sums[11][41] , \sums[11][40] , \sums[11][39] , 
    \sums[11][38] , \sums[11][37] , \sums[11][36] , \sums[11][35] , \sums[11][34] , 
    \sums[11][33] , \sums[11][32] , \sums[11][31] , \sums[11][30] , \sums[11][29] , 
    \sums[11][28] , \sums[11][27] , \sums[11][26] , \sums[11][25] , \sums[11][24] , 
    \sums[11][23] , \sums[11][22] , \sums[11][21] , \sums[11][20] , \sums[11][19] , 
    \sums[11][18] , \sums[11][17] , \sums[11][16] , \sums[11][15] , \sums[11][14] , 
    \sums[11][13] , \sums[11][12] , \sums[11][11] , \sums[11][10] , \sums[11][9] , 
    \sums[11][8] , \sums[11][7] , \sums[11][6] , n_2_0, uc_2184, uc_2185, uc_2186, 
    uc_2187, uc_2188}));
CSA__0_72 CSA18 (.u ({\sums[18][63] , \sums[18][62] , \sums[18][61] , \sums[18][60] , 
    \sums[18][59] , \sums[18][58] , \sums[18][57] , \sums[18][56] , \sums[18][55] , 
    \sums[18][54] , \sums[18][53] , \sums[18][52] , \sums[18][51] , \sums[18][50] , 
    \sums[18][49] , \sums[18][48] , \sums[18][47] , \sums[18][46] , \sums[18][45] , 
    \sums[18][44] , \sums[18][43] , \sums[18][42] , \sums[18][41] , \sums[18][40] , 
    \sums[18][39] , \sums[18][38] , \sums[18][37] , \sums[18][36] , \sums[18][35] , 
    \sums[18][34] , \sums[18][33] , \sums[18][32] , \sums[18][31] , \sums[18][30] , 
    \sums[18][29] , \sums[18][28] , \sums[18][27] , \sums[18][26] , \sums[18][25] , 
    \sums[18][24] , \sums[18][23] , \sums[18][22] , \sums[18][21] , \sums[18][20] , 
    \sums[18][19] , \sums[18][18] , \sums[18][17] , \sums[18][16] , \sums[18][15] , 
    \sums[18][14] , \sums[18][13] , \sums[18][12] , \sums[18][11] , \sums[18][10] , 
    \sums[18][9] , uc_2106, uc_2107, uc_2108, uc_2109, uc_2110, uc_2111, uc_2112, 
    uc_2113, uc_2114}), .v ({\couts[18][63] , \couts[18][62] , \couts[18][61] , \couts[18][60] , 
    \couts[18][59] , \couts[18][58] , \couts[18][57] , \couts[18][56] , \couts[18][55] , 
    \couts[18][54] , \couts[18][53] , \couts[18][52] , \couts[18][51] , \couts[18][50] , 
    \couts[18][49] , \couts[18][48] , \couts[18][47] , \couts[18][46] , \couts[18][45] , 
    \couts[18][44] , \couts[18][43] , \couts[18][42] , \couts[18][41] , \couts[18][40] , 
    \couts[18][39] , \couts[18][38] , \couts[18][37] , \couts[18][36] , \couts[18][35] , 
    \couts[18][34] , \couts[18][33] , \couts[18][32] , \couts[18][31] , \couts[18][30] , 
    \couts[18][29] , \couts[18][28] , \couts[18][27] , \couts[18][26] , \couts[18][25] , 
    \couts[18][24] , \couts[18][23] , \couts[18][22] , \couts[18][21] , \couts[18][20] , 
    \couts[18][19] , \couts[18][18] , \couts[18][17] , \couts[18][16] , \couts[18][15] , 
    \couts[18][14] , \couts[18][13] , \couts[18][12] , \couts[18][11] , \couts[18][10] , 
    uc_2115, uc_2116, uc_2117, uc_2118, uc_2119, uc_2120, uc_2121, uc_2122, uc_2123, 
    uc_2124}), .x ({\couts[11][63] , \couts[11][62] , \couts[11][61] , \couts[11][60] , 
    \couts[11][59] , \couts[11][58] , \couts[11][57] , \couts[11][56] , \couts[11][55] , 
    \couts[11][54] , \couts[11][53] , \couts[11][52] , \couts[11][51] , \couts[11][50] , 
    \couts[11][49] , \couts[11][48] , \couts[11][47] , \couts[11][46] , \couts[11][45] , 
    \couts[11][44] , \couts[11][43] , \couts[11][42] , \couts[11][41] , \couts[11][40] , 
    \couts[11][39] , \couts[11][38] , \couts[11][37] , \couts[11][36] , \couts[11][35] , 
    \couts[11][34] , \couts[11][33] , \couts[11][32] , \couts[11][31] , \couts[11][30] , 
    \couts[11][29] , \couts[11][28] , \couts[11][27] , \couts[11][26] , \couts[11][25] , 
    \couts[11][24] , \couts[11][23] , \couts[11][22] , \couts[11][21] , \couts[11][20] , 
    \couts[11][19] , \couts[11][18] , \couts[11][17] , \couts[11][16] , \couts[11][15] , 
    \couts[11][14] , \couts[11][13] , \couts[11][12] , \couts[11][11] , \couts[11][10] , 
    \couts[11][9] , uc_2041, uc_2042, uc_2043, uc_2044, uc_2045, uc_2046, uc_2047, 
    uc_2048, uc_2049}), .y ({\sums[12][63] , uc_2050, uc_2051, uc_2052, uc_2053, 
    uc_2054, uc_2055, uc_2056, uc_2057, uc_2058, uc_2059, uc_2060, uc_2061, uc_2062, 
    uc_2063, uc_2064, uc_2065, uc_2066, uc_2067, \sums[12][44] , \sums[12][43] , 
    \sums[12][42] , \sums[12][41] , \sums[12][40] , \sums[12][39] , \sums[12][38] , 
    \sums[12][37] , \sums[12][36] , \sums[12][35] , \sums[12][34] , \sums[12][33] , 
    \sums[12][32] , \sums[12][31] , \sums[12][30] , \sums[12][29] , \sums[12][28] , 
    \sums[12][27] , \sums[12][26] , \sums[12][25] , \sums[12][24] , \sums[12][23] , 
    \sums[12][22] , \sums[12][21] , \sums[12][20] , \sums[12][19] , \sums[12][18] , 
    \sums[12][17] , \sums[12][16] , \sums[12][15] , \sums[12][14] , \sums[12][13] , 
    \sums[12][12] , \sums[12][11] , \sums[3][10] , \pp[9][9] , uc_2068, uc_2069, 
    uc_2070, uc_2071, uc_2072, uc_2073, uc_2074, uc_2075, uc_2076}), .z ({\couts[12][63] , 
    uc_2077, uc_2078, uc_2079, uc_2080, uc_2081, uc_2082, uc_2083, uc_2084, uc_2085, 
    uc_2086, uc_2087, uc_2088, uc_2089, uc_2090, uc_2091, uc_2092, uc_2093, \couts[12][45] , 
    \couts[12][44] , \couts[12][43] , \couts[12][42] , \couts[12][41] , \couts[12][40] , 
    \couts[12][39] , \couts[12][38] , \couts[12][37] , \couts[12][36] , \couts[12][35] , 
    \couts[12][34] , \couts[12][33] , \couts[12][32] , \couts[12][31] , \couts[12][30] , 
    \couts[12][29] , \couts[12][28] , \couts[12][27] , \couts[12][26] , \couts[12][25] , 
    \couts[12][24] , \couts[12][23] , \couts[12][22] , \couts[12][21] , \couts[12][20] , 
    \couts[12][19] , \couts[12][18] , \couts[12][17] , \couts[12][16] , \couts[12][15] , 
    \couts[12][14] , \couts[12][13] , \couts[12][12] , uc_2094, uc_2095, uc_2096, 
    uc_2097, uc_2098, uc_2099, uc_2100, uc_2101, uc_2102, uc_2103, uc_2104, uc_2105}));
CSA__2_11 CSA3 (.u ({\sums[3][63] , uc_1979, uc_1980, uc_1981, uc_1982, uc_1983, 
    uc_1984, uc_1985, uc_1986, uc_1987, uc_1988, uc_1989, uc_1990, uc_1991, uc_1992, 
    uc_1993, uc_1994, uc_1995, uc_1996, uc_1997, uc_1998, uc_1999, \sums[3][41] , 
    \sums[3][40] , \sums[3][39] , \sums[3][38] , \sums[3][37] , \sums[3][36] , \sums[3][35] , 
    \sums[3][34] , \sums[3][33] , \sums[3][32] , \sums[3][31] , \sums[3][30] , \sums[3][29] , 
    \sums[3][28] , \sums[3][27] , \sums[3][26] , \sums[3][25] , \sums[3][24] , \sums[3][23] , 
    \sums[3][22] , \sums[3][21] , \sums[3][20] , \sums[3][19] , \sums[3][18] , \sums[3][17] , 
    \sums[3][16] , \sums[3][15] , \sums[3][14] , \sums[3][13] , \sums[3][12] , \sums[3][11] , 
    \sums[3][10] , uc_2000, uc_2001, uc_2002, uc_2003, uc_2004, uc_2005, uc_2006, 
    uc_2007, uc_2008, uc_2009}), .v ({\couts[3][63] , uc_2010, uc_2011, uc_2012, 
    uc_2013, uc_2014, uc_2015, uc_2016, uc_2017, uc_2018, uc_2019, uc_2020, uc_2021, 
    uc_2022, uc_2023, uc_2024, uc_2025, uc_2026, uc_2027, uc_2028, uc_2029, \couts[3][42] , 
    \couts[3][41] , \couts[3][40] , \couts[3][39] , \couts[3][38] , \couts[3][37] , 
    \couts[3][36] , \couts[3][35] , \couts[3][34] , \couts[3][33] , \couts[3][32] , 
    \couts[3][31] , \couts[3][30] , \couts[3][29] , \couts[3][28] , \couts[3][27] , 
    \couts[3][26] , \couts[3][25] , \couts[3][24] , \couts[3][23] , \couts[3][22] , 
    \couts[3][21] , \couts[3][20] , \couts[3][19] , \couts[3][18] , \couts[3][17] , 
    \couts[3][16] , \couts[3][15] , \couts[3][14] , \couts[3][13] , \couts[3][12] , 
    \couts[3][11] , uc_2030, uc_2031, uc_2032, uc_2033, uc_2034, uc_2035, uc_2036, 
    uc_2037, uc_2038, uc_2039, uc_2040}), .x ({uc_1882, \pp[9][63] , uc_1883, uc_1884, 
    uc_1885, uc_1886, uc_1887, uc_1888, uc_1889, uc_1890, uc_1891, uc_1892, uc_1893, 
    uc_1894, uc_1895, uc_1896, uc_1897, uc_1898, uc_1899, uc_1900, uc_1901, uc_1902, 
    uc_1903, uc_1904, \pp[9][39] , \pp[9][38] , \pp[9][37] , \pp[9][36] , \pp[9][35] , 
    \pp[9][34] , \pp[9][33] , \pp[9][32] , \pp[9][31] , \pp[9][30] , \pp[9][29] , 
    \pp[9][28] , \pp[9][27] , \pp[9][26] , \pp[9][25] , \pp[9][24] , \pp[9][23] , 
    \pp[9][22] , \pp[9][21] , \pp[9][20] , \pp[9][19] , \pp[9][18] , \pp[9][17] , 
    \pp[9][16] , \pp[9][15] , \pp[9][14] , \pp[9][13] , \pp[9][12] , \pp[9][11] , 
    \pp[9][10] , uc_1905, uc_1906, uc_1907, uc_1908, uc_1909, uc_1910, uc_1911, uc_1912, 
    uc_1913, uc_1914}), .y ({uc_1915, \pp[10][63] , uc_1916, uc_1917, uc_1918, uc_1919, 
    uc_1920, uc_1921, uc_1922, uc_1923, uc_1924, uc_1925, uc_1926, uc_1927, uc_1928, 
    uc_1929, uc_1930, uc_1931, uc_1932, uc_1933, uc_1934, uc_1935, uc_1936, \pp[10][40] , 
    \pp[10][39] , \pp[10][38] , \pp[10][37] , \pp[10][36] , \pp[10][35] , \pp[10][34] , 
    \pp[10][33] , \pp[10][32] , \pp[10][31] , \pp[10][30] , \pp[10][29] , \pp[10][28] , 
    \pp[10][27] , \pp[10][26] , \pp[10][25] , \pp[10][24] , \pp[10][23] , \pp[10][22] , 
    \pp[10][21] , \pp[10][20] , \pp[10][19] , \pp[10][18] , \pp[10][17] , \pp[10][16] , 
    \pp[10][15] , \pp[10][14] , \pp[10][13] , \pp[10][12] , \pp[10][11] , \pp[10][10] , 
    uc_1937, uc_1938, uc_1939, uc_1940, uc_1941, uc_1942, uc_1943, uc_1944, uc_1945, 
    uc_1946}), .z ({uc_1947, \pp[11][63] , uc_1948, uc_1949, uc_1950, uc_1951, uc_1952, 
    uc_1953, uc_1954, uc_1955, uc_1956, uc_1957, uc_1958, uc_1959, uc_1960, uc_1961, 
    uc_1962, uc_1963, uc_1964, uc_1965, uc_1966, uc_1967, \pp[11][41] , \pp[11][40] , 
    \pp[11][39] , \pp[11][38] , \pp[11][37] , \pp[11][36] , \pp[11][35] , \pp[11][34] , 
    \pp[11][33] , \pp[11][32] , \pp[11][31] , \pp[11][30] , \pp[11][29] , \pp[11][28] , 
    \pp[11][27] , \pp[11][26] , \pp[11][25] , \pp[11][24] , \pp[11][23] , \pp[11][22] , 
    \pp[11][21] , \pp[11][20] , \pp[11][19] , \pp[11][18] , \pp[11][17] , \pp[11][16] , 
    \pp[11][15] , \pp[11][14] , \pp[11][13] , \pp[11][12] , \pp[11][11] , uc_1968, 
    uc_1969, uc_1970, uc_1971, uc_1972, uc_1973, uc_1974, uc_1975, uc_1976, uc_1977, 
    uc_1978}));
CSA__2_8 CSA12 (.u ({\sums[12][63] , uc_1824, uc_1825, uc_1826, uc_1827, uc_1828, 
    uc_1829, uc_1830, uc_1831, uc_1832, uc_1833, uc_1834, uc_1835, uc_1836, uc_1837, 
    uc_1838, uc_1839, uc_1840, uc_1841, \sums[12][44] , \sums[12][43] , \sums[12][42] , 
    \sums[12][41] , \sums[12][40] , \sums[12][39] , \sums[12][38] , \sums[12][37] , 
    \sums[12][36] , \sums[12][35] , \sums[12][34] , \sums[12][33] , \sums[12][32] , 
    \sums[12][31] , \sums[12][30] , \sums[12][29] , \sums[12][28] , \sums[12][27] , 
    \sums[12][26] , \sums[12][25] , \sums[12][24] , \sums[12][23] , \sums[12][22] , 
    \sums[12][21] , \sums[12][20] , \sums[12][19] , \sums[12][18] , \sums[12][17] , 
    \sums[12][16] , \sums[12][15] , \sums[12][14] , \sums[12][13] , \sums[12][12] , 
    \sums[12][11] , uc_1842, uc_1843, uc_1844, uc_1845, uc_1846, uc_1847, uc_1848, 
    uc_1849, uc_1850, uc_1851, uc_1852}), .v ({\couts[12][63] , uc_1853, uc_1854, 
    uc_1855, uc_1856, uc_1857, uc_1858, uc_1859, uc_1860, uc_1861, uc_1862, uc_1863, 
    uc_1864, uc_1865, uc_1866, uc_1867, uc_1868, uc_1869, \couts[12][45] , \couts[12][44] , 
    \couts[12][43] , \couts[12][42] , \couts[12][41] , \couts[12][40] , \couts[12][39] , 
    \couts[12][38] , \couts[12][37] , \couts[12][36] , \couts[12][35] , \couts[12][34] , 
    \couts[12][33] , \couts[12][32] , \couts[12][31] , \couts[12][30] , \couts[12][29] , 
    \couts[12][28] , \couts[12][27] , \couts[12][26] , \couts[12][25] , \couts[12][24] , 
    \couts[12][23] , \couts[12][22] , \couts[12][21] , \couts[12][20] , \couts[12][19] , 
    \couts[12][18] , \couts[12][17] , \couts[12][16] , \couts[12][15] , \couts[12][14] , 
    \couts[12][13] , \couts[12][12] , uc_1870, uc_1871, uc_1872, uc_1873, uc_1874, 
    uc_1875, uc_1876, uc_1877, uc_1878, uc_1879, uc_1880, uc_1881}), .x ({\sums[3][63] , 
    uc_1731, uc_1732, uc_1733, uc_1734, uc_1735, uc_1736, uc_1737, uc_1738, uc_1739, 
    uc_1740, uc_1741, uc_1742, uc_1743, uc_1744, uc_1745, uc_1746, uc_1747, uc_1748, 
    uc_1749, uc_1750, uc_1751, \sums[3][41] , \sums[3][40] , \sums[3][39] , \sums[3][38] , 
    \sums[3][37] , \sums[3][36] , \sums[3][35] , \sums[3][34] , \sums[3][33] , \sums[3][32] , 
    \sums[3][31] , \sums[3][30] , \sums[3][29] , \sums[3][28] , \sums[3][27] , \sums[3][26] , 
    \sums[3][25] , \sums[3][24] , \sums[3][23] , \sums[3][22] , \sums[3][21] , \sums[3][20] , 
    \sums[3][19] , \sums[3][18] , \sums[3][17] , \sums[3][16] , \sums[3][15] , \sums[3][14] , 
    \sums[3][13] , \sums[3][12] , \sums[3][11] , uc_1752, uc_1753, uc_1754, uc_1755, 
    uc_1756, uc_1757, uc_1758, uc_1759, uc_1760, uc_1761, uc_1762}), .y ({\couts[3][63] , 
    uc_1763, uc_1764, uc_1765, uc_1766, uc_1767, uc_1768, uc_1769, uc_1770, uc_1771, 
    uc_1772, uc_1773, uc_1774, uc_1775, uc_1776, uc_1777, uc_1778, uc_1779, uc_1780, 
    uc_1781, uc_1782, \couts[3][42] , \couts[3][41] , \couts[3][40] , \couts[3][39] , 
    \couts[3][38] , \couts[3][37] , \couts[3][36] , \couts[3][35] , \couts[3][34] , 
    \couts[3][33] , \couts[3][32] , \couts[3][31] , \couts[3][30] , \couts[3][29] , 
    \couts[3][28] , \couts[3][27] , \couts[3][26] , \couts[3][25] , \couts[3][24] , 
    \couts[3][23] , \couts[3][22] , \couts[3][21] , \couts[3][20] , \couts[3][19] , 
    \couts[3][18] , \couts[3][17] , \couts[3][16] , \couts[3][15] , \couts[3][14] , 
    \couts[3][13] , \couts[3][12] , \couts[3][11] , uc_1783, uc_1784, uc_1785, uc_1786, 
    uc_1787, uc_1788, uc_1789, uc_1790, uc_1791, uc_1792, uc_1793}), .z ({\sums[4][63] , 
    uc_1794, uc_1795, uc_1796, uc_1797, uc_1798, uc_1799, uc_1800, uc_1801, uc_1802, 
    uc_1803, uc_1804, uc_1805, uc_1806, uc_1807, uc_1808, uc_1809, uc_1810, uc_1811, 
    \sums[4][44] , \sums[4][43] , \sums[4][42] , \sums[4][41] , \sums[4][40] , \sums[4][39] , 
    \sums[4][38] , \sums[4][37] , \sums[4][36] , \sums[4][35] , \sums[4][34] , \sums[4][33] , 
    \sums[4][32] , \sums[4][31] , \sums[4][30] , \sums[4][29] , \sums[4][28] , \sums[4][27] , 
    \sums[4][26] , \sums[4][25] , \sums[4][24] , \sums[4][23] , \sums[4][22] , \sums[4][21] , 
    \sums[4][20] , \sums[4][19] , \sums[4][18] , \sums[4][17] , \sums[4][16] , \sums[4][15] , 
    \sums[4][14] , \sums[4][13] , \sums[4][12] , uc_1812, uc_1813, uc_1814, uc_1815, 
    uc_1816, uc_1817, uc_1818, uc_1819, uc_1820, uc_1821, uc_1822, uc_1823}));
CSA__2_5 CSA11 (.u ({\sums[11][63] , \sums[11][62] , \sums[11][61] , \sums[11][60] , 
    \sums[11][59] , \sums[11][58] , \sums[11][57] , \sums[11][56] , \sums[11][55] , 
    \sums[11][54] , \sums[11][53] , \sums[11][52] , \sums[11][51] , \sums[11][50] , 
    \sums[11][49] , \sums[11][48] , \sums[11][47] , \sums[11][46] , \sums[11][45] , 
    \sums[11][44] , \sums[11][43] , \sums[11][42] , \sums[11][41] , \sums[11][40] , 
    \sums[11][39] , \sums[11][38] , \sums[11][37] , \sums[11][36] , \sums[11][35] , 
    \sums[11][34] , \sums[11][33] , \sums[11][32] , \sums[11][31] , \sums[11][30] , 
    \sums[11][29] , \sums[11][28] , \sums[11][27] , \sums[11][26] , \sums[11][25] , 
    \sums[11][24] , \sums[11][23] , \sums[11][22] , \sums[11][21] , \sums[11][20] , 
    \sums[11][19] , \sums[11][18] , \sums[11][17] , \sums[11][16] , \sums[11][15] , 
    \sums[11][14] , \sums[11][13] , \sums[11][12] , \sums[11][11] , \sums[11][10] , 
    \sums[11][9] , \sums[11][8] , \sums[11][7] , \sums[11][6] , uc_1718, uc_1719, 
    uc_1720, uc_1721, uc_1722, uc_1723}), .v ({\couts[11][63] , \couts[11][62] , 
    \couts[11][61] , \couts[11][60] , \couts[11][59] , \couts[11][58] , \couts[11][57] , 
    \couts[11][56] , \couts[11][55] , \couts[11][54] , \couts[11][53] , \couts[11][52] , 
    \couts[11][51] , \couts[11][50] , \couts[11][49] , \couts[11][48] , \couts[11][47] , 
    \couts[11][46] , \couts[11][45] , \couts[11][44] , \couts[11][43] , \couts[11][42] , 
    \couts[11][41] , \couts[11][40] , \couts[11][39] , \couts[11][38] , \couts[11][37] , 
    \couts[11][36] , \couts[11][35] , \couts[11][34] , \couts[11][33] , \couts[11][32] , 
    \couts[11][31] , \couts[11][30] , \couts[11][29] , \couts[11][28] , \couts[11][27] , 
    \couts[11][26] , \couts[11][25] , \couts[11][24] , \couts[11][23] , \couts[11][22] , 
    \couts[11][21] , \couts[11][20] , \couts[11][19] , \couts[11][18] , \couts[11][17] , 
    \couts[11][16] , \couts[11][15] , \couts[11][14] , \couts[11][13] , \couts[11][12] , 
    \couts[11][11] , \couts[11][10] , \couts[11][9] , \sums[18][8] , \sums[18][7] , 
    uc_1724, uc_1725, uc_1726, uc_1727, uc_1728, uc_1729, uc_1730}), .x ({\couts[1][37] , 
    \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , 
    \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , 
    \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , 
    \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , 
    \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , \couts[1][37] , 
    \couts[1][37] , \couts[1][36] , \couts[1][35] , \couts[1][34] , \couts[1][33] , 
    \couts[1][32] , \couts[1][31] , \couts[1][30] , \couts[1][29] , \couts[1][28] , 
    \couts[1][27] , \couts[1][26] , \couts[1][25] , \couts[1][24] , \couts[1][23] , 
    \couts[1][22] , \couts[1][21] , \couts[1][20] , \couts[1][19] , \couts[1][18] , 
    \couts[1][17] , \couts[1][16] , \couts[1][15] , \couts[1][14] , \couts[1][13] , 
    \couts[1][12] , \couts[1][11] , \couts[1][10] , \couts[1][9] , \couts[1][8] , 
    \couts[1][7] , \couts[1][6] , uc_1651, uc_1652, uc_1653, uc_1654, uc_1655, uc_1656})
    , .y ({\sums[2][63] , uc_1657, uc_1658, uc_1659, uc_1660, uc_1661, uc_1662, uc_1663, 
    uc_1664, uc_1665, uc_1666, uc_1667, uc_1668, uc_1669, uc_1670, uc_1671, uc_1672, 
    uc_1673, uc_1674, uc_1675, uc_1676, uc_1677, uc_1678, uc_1679, uc_1680, \sums[2][38] , 
    \sums[2][37] , \sums[2][36] , \sums[2][35] , \sums[2][34] , \sums[2][33] , \sums[2][32] , 
    \sums[2][31] , \sums[2][30] , \sums[2][29] , \sums[2][28] , \sums[2][27] , \sums[2][26] , 
    \sums[2][25] , \sums[2][24] , \sums[2][23] , \sums[2][22] , \sums[2][21] , \sums[2][20] , 
    \sums[2][19] , \sums[2][18] , \sums[2][17] , \sums[2][16] , \sums[2][15] , \sums[2][14] , 
    \sums[2][13] , \sums[2][12] , \sums[2][11] , \sums[2][10] , \sums[2][9] , \sums[2][8] , 
    \sums[2][7] , \pp[6][6] , uc_1681, uc_1682, uc_1683, uc_1684, uc_1685, uc_1686})
    , .z ({\couts[2][63] , uc_1687, uc_1688, uc_1689, uc_1690, uc_1691, uc_1692, 
    uc_1693, uc_1694, uc_1695, uc_1696, uc_1697, uc_1698, uc_1699, uc_1700, uc_1701, 
    uc_1702, uc_1703, uc_1704, uc_1705, uc_1706, uc_1707, uc_1708, uc_1709, \couts[2][39] , 
    \couts[2][38] , \couts[2][37] , \couts[2][36] , \couts[2][35] , \couts[2][34] , 
    \couts[2][33] , \couts[2][32] , \couts[2][31] , \couts[2][30] , \couts[2][29] , 
    \couts[2][28] , \couts[2][27] , \couts[2][26] , \couts[2][25] , \couts[2][24] , 
    \couts[2][23] , \couts[2][22] , \couts[2][21] , \couts[2][20] , \couts[2][19] , 
    \couts[2][18] , \couts[2][17] , \couts[2][16] , \couts[2][15] , \couts[2][14] , 
    \couts[2][13] , \couts[2][12] , \couts[2][11] , \couts[2][10] , \couts[2][9] , 
    \couts[2][8] , uc_1710, uc_1711, uc_1712, uc_1713, uc_1714, uc_1715, uc_1716, 
    uc_1717}));
CSA__2_2 CSA2 (.u ({\sums[2][63] , uc_1589, uc_1590, uc_1591, uc_1592, uc_1593, uc_1594, 
    uc_1595, uc_1596, uc_1597, uc_1598, uc_1599, uc_1600, uc_1601, uc_1602, uc_1603, 
    uc_1604, uc_1605, uc_1606, uc_1607, uc_1608, uc_1609, uc_1610, uc_1611, uc_1612, 
    \sums[2][38] , \sums[2][37] , \sums[2][36] , \sums[2][35] , \sums[2][34] , \sums[2][33] , 
    \sums[2][32] , \sums[2][31] , \sums[2][30] , \sums[2][29] , \sums[2][28] , \sums[2][27] , 
    \sums[2][26] , \sums[2][25] , \sums[2][24] , \sums[2][23] , \sums[2][22] , \sums[2][21] , 
    \sums[2][20] , \sums[2][19] , \sums[2][18] , \sums[2][17] , \sums[2][16] , \sums[2][15] , 
    \sums[2][14] , \sums[2][13] , \sums[2][12] , \sums[2][11] , \sums[2][10] , \sums[2][9] , 
    \sums[2][8] , \sums[2][7] , uc_1613, uc_1614, uc_1615, uc_1616, uc_1617, uc_1618, 
    uc_1619}), .v ({\couts[2][63] , uc_1620, uc_1621, uc_1622, uc_1623, uc_1624, 
    uc_1625, uc_1626, uc_1627, uc_1628, uc_1629, uc_1630, uc_1631, uc_1632, uc_1633, 
    uc_1634, uc_1635, uc_1636, uc_1637, uc_1638, uc_1639, uc_1640, uc_1641, uc_1642, 
    \couts[2][39] , \couts[2][38] , \couts[2][37] , \couts[2][36] , \couts[2][35] , 
    \couts[2][34] , \couts[2][33] , \couts[2][32] , \couts[2][31] , \couts[2][30] , 
    \couts[2][29] , \couts[2][28] , \couts[2][27] , \couts[2][26] , \couts[2][25] , 
    \couts[2][24] , \couts[2][23] , \couts[2][22] , \couts[2][21] , \couts[2][20] , 
    \couts[2][19] , \couts[2][18] , \couts[2][17] , \couts[2][16] , \couts[2][15] , 
    \couts[2][14] , \couts[2][13] , \couts[2][12] , \couts[2][11] , \couts[2][10] , 
    \couts[2][9] , \couts[2][8] , uc_1643, uc_1644, uc_1645, uc_1646, uc_1647, uc_1648, 
    uc_1649, uc_1650}), .x ({\pp[6][63] , uc_1492, uc_1493, uc_1494, uc_1495, uc_1496, 
    uc_1497, uc_1498, uc_1499, uc_1500, uc_1501, uc_1502, uc_1503, uc_1504, uc_1505, 
    uc_1506, uc_1507, uc_1508, uc_1509, uc_1510, uc_1511, uc_1512, uc_1513, uc_1514, 
    uc_1515, uc_1516, uc_1517, \pp[6][36] , \pp[6][35] , \pp[6][34] , \pp[6][33] , 
    \pp[6][32] , \pp[6][31] , \pp[6][30] , \pp[6][29] , \pp[6][28] , \pp[6][27] , 
    \pp[6][26] , \pp[6][25] , \pp[6][24] , \pp[6][23] , \pp[6][22] , \pp[6][21] , 
    \pp[6][20] , \pp[6][19] , \pp[6][18] , \pp[6][17] , \pp[6][16] , \pp[6][15] , 
    \pp[6][14] , \pp[6][13] , \pp[6][12] , \pp[6][11] , \pp[6][10] , \pp[6][9] , 
    \pp[6][8] , \pp[6][7] , uc_1518, uc_1519, uc_1520, uc_1521, uc_1522, uc_1523, 
    uc_1524}), .y ({\pp[7][63] , uc_1525, uc_1526, uc_1527, uc_1528, uc_1529, uc_1530, 
    uc_1531, uc_1532, uc_1533, uc_1534, uc_1535, uc_1536, uc_1537, uc_1538, uc_1539, 
    uc_1540, uc_1541, uc_1542, uc_1543, uc_1544, uc_1545, uc_1546, uc_1547, uc_1548, 
    uc_1549, \pp[7][37] , \pp[7][36] , \pp[7][35] , \pp[7][34] , \pp[7][33] , \pp[7][32] , 
    \pp[7][31] , \pp[7][30] , \pp[7][29] , \pp[7][28] , \pp[7][27] , \pp[7][26] , 
    \pp[7][25] , \pp[7][24] , \pp[7][23] , \pp[7][22] , \pp[7][21] , \pp[7][20] , 
    \pp[7][19] , \pp[7][18] , \pp[7][17] , \pp[7][16] , \pp[7][15] , \pp[7][14] , 
    \pp[7][13] , \pp[7][12] , \pp[7][11] , \pp[7][10] , \pp[7][9] , \pp[7][8] , \pp[7][7] , 
    uc_1550, uc_1551, uc_1552, uc_1553, uc_1554, uc_1555, uc_1556}), .z ({\pp[8][63] , 
    uc_1557, uc_1558, uc_1559, uc_1560, uc_1561, uc_1562, uc_1563, uc_1564, uc_1565, 
    uc_1566, uc_1567, uc_1568, uc_1569, uc_1570, uc_1571, uc_1572, uc_1573, uc_1574, 
    uc_1575, uc_1576, uc_1577, uc_1578, uc_1579, uc_1580, \pp[8][38] , \pp[8][37] , 
    \pp[8][36] , \pp[8][35] , \pp[8][34] , \pp[8][33] , \pp[8][32] , \pp[8][31] , 
    \pp[8][30] , \pp[8][29] , \pp[8][28] , \pp[8][27] , \pp[8][26] , \pp[8][25] , 
    \pp[8][24] , \pp[8][23] , \pp[8][22] , \pp[8][21] , \pp[8][20] , \pp[8][19] , 
    \pp[8][18] , \pp[8][17] , \pp[8][16] , \pp[8][15] , \pp[8][14] , \pp[8][13] , 
    \pp[8][12] , \pp[8][11] , \pp[8][10] , \pp[8][9] , \pp[8][8] , uc_1581, uc_1582, 
    uc_1583, uc_1584, uc_1585, uc_1586, uc_1587, uc_1588}));
CSA__0_69 CSA4 (.u ({\sums[4][63] , uc_1430, uc_1431, uc_1432, uc_1433, uc_1434, 
    uc_1435, uc_1436, uc_1437, uc_1438, uc_1439, uc_1440, uc_1441, uc_1442, uc_1443, 
    uc_1444, uc_1445, uc_1446, uc_1447, \sums[4][44] , \sums[4][43] , \sums[4][42] , 
    \sums[4][41] , \sums[4][40] , \sums[4][39] , \sums[4][38] , \sums[4][37] , \sums[4][36] , 
    \sums[4][35] , \sums[4][34] , \sums[4][33] , \sums[4][32] , \sums[4][31] , \sums[4][30] , 
    \sums[4][29] , \sums[4][28] , \sums[4][27] , \sums[4][26] , \sums[4][25] , \sums[4][24] , 
    \sums[4][23] , \sums[4][22] , \sums[4][21] , \sums[4][20] , \sums[4][19] , \sums[4][18] , 
    \sums[4][17] , \sums[4][16] , \sums[4][15] , \sums[4][14] , \sums[4][13] , uc_1448, 
    uc_1449, uc_1450, uc_1451, uc_1452, uc_1453, uc_1454, uc_1455, uc_1456, uc_1457, 
    uc_1458, uc_1459, uc_1460}), .v ({\couts[4][63] , uc_1461, uc_1462, uc_1463, 
    uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, uc_1469, uc_1470, uc_1471, uc_1472, 
    uc_1473, uc_1474, uc_1475, uc_1476, uc_1477, \couts[4][45] , \couts[4][44] , 
    \couts[4][43] , \couts[4][42] , \couts[4][41] , \couts[4][40] , \couts[4][39] , 
    \couts[4][38] , \couts[4][37] , \couts[4][36] , \couts[4][35] , \couts[4][34] , 
    \couts[4][33] , \couts[4][32] , \couts[4][31] , \couts[4][30] , \couts[4][29] , 
    \couts[4][28] , \couts[4][27] , \couts[4][26] , \couts[4][25] , \couts[4][24] , 
    \couts[4][23] , \couts[4][22] , \couts[4][21] , \couts[4][20] , \couts[4][19] , 
    \couts[4][18] , \couts[4][17] , \couts[4][16] , \couts[4][15] , \sums[13][14] , 
    uc_1478, uc_1479, uc_1480, uc_1481, uc_1482, uc_1483, uc_1484, uc_1485, uc_1486, 
    uc_1487, uc_1488, uc_1489, uc_1490, uc_1491}), .x ({uc_1333, \pp[12][62] , uc_1334, 
    uc_1335, uc_1336, uc_1337, uc_1338, uc_1339, uc_1340, uc_1341, uc_1342, uc_1343, 
    uc_1344, uc_1345, uc_1346, uc_1347, uc_1348, uc_1349, uc_1350, uc_1351, uc_1352, 
    \pp[12][42] , \pp[12][41] , \pp[12][40] , \pp[12][39] , \pp[12][38] , \pp[12][37] , 
    \pp[12][36] , \pp[12][35] , \pp[12][34] , \pp[12][33] , \pp[12][32] , \pp[12][31] , 
    \pp[12][30] , \pp[12][29] , \pp[12][28] , \pp[12][27] , \pp[12][26] , \pp[12][25] , 
    \pp[12][24] , \pp[12][23] , \pp[12][22] , \pp[12][21] , \pp[12][20] , \pp[12][19] , 
    \pp[12][18] , \pp[12][17] , \pp[12][16] , \pp[12][15] , \pp[12][14] , \pp[12][13] , 
    uc_1353, uc_1354, uc_1355, uc_1356, uc_1357, uc_1358, uc_1359, uc_1360, uc_1361, 
    uc_1362, uc_1363, uc_1364, uc_1365}), .y ({uc_1366, \pp[13][62] , uc_1367, uc_1368, 
    uc_1369, uc_1370, uc_1371, uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, uc_1377, 
    uc_1378, uc_1379, uc_1380, uc_1381, uc_1382, uc_1383, uc_1384, \pp[13][43] , 
    \pp[13][42] , \pp[13][41] , \pp[13][40] , \pp[13][39] , \pp[13][38] , \pp[13][37] , 
    \pp[13][36] , \pp[13][35] , \pp[13][34] , \pp[13][33] , \pp[13][32] , \pp[13][31] , 
    \pp[13][30] , \pp[13][29] , \pp[13][28] , \pp[13][27] , \pp[13][26] , \pp[13][25] , 
    \pp[13][24] , \pp[13][23] , \pp[13][22] , \pp[13][21] , \pp[13][20] , \pp[13][19] , 
    \pp[13][18] , \pp[13][17] , \pp[13][16] , \pp[13][15] , \pp[13][14] , \pp[13][13] , 
    uc_1385, uc_1386, uc_1387, uc_1388, uc_1389, uc_1390, uc_1391, uc_1392, uc_1393, 
    uc_1394, uc_1395, uc_1396, uc_1397}), .z ({uc_1398, \pp[14][62] , uc_1399, uc_1400, 
    uc_1401, uc_1402, uc_1403, uc_1404, uc_1405, uc_1406, uc_1407, uc_1408, uc_1409, 
    uc_1410, uc_1411, uc_1412, uc_1413, uc_1414, uc_1415, \pp[14][44] , \pp[14][43] , 
    \pp[14][42] , \pp[14][41] , \pp[14][40] , \pp[14][39] , \pp[14][38] , \pp[14][37] , 
    \pp[14][36] , \pp[14][35] , \pp[14][34] , \pp[14][33] , \pp[14][32] , \pp[14][31] , 
    \pp[14][30] , \pp[14][29] , \pp[14][28] , \pp[14][27] , \pp[14][26] , \pp[14][25] , 
    \pp[14][24] , \pp[14][23] , \pp[14][22] , \pp[14][21] , \pp[14][20] , \pp[14][19] , 
    \pp[14][18] , \pp[14][17] , \pp[14][16] , \pp[14][15] , \pp[14][14] , uc_1416, 
    uc_1417, uc_1418, uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, uc_1424, uc_1425, 
    uc_1426, uc_1427, uc_1428, uc_1429}));
CSA__1_5 CSA5 (.u ({\sums[5][63] , uc_1271, uc_1272, uc_1273, uc_1274, uc_1275, uc_1276, 
    uc_1277, uc_1278, uc_1279, uc_1280, uc_1281, uc_1282, uc_1283, uc_1284, uc_1285, 
    \sums[5][47] , \sums[5][46] , \sums[5][45] , \sums[5][44] , \sums[5][43] , \sums[5][42] , 
    \sums[5][41] , \sums[5][40] , \sums[5][39] , \sums[5][38] , \sums[5][37] , \sums[5][36] , 
    \sums[5][35] , \sums[5][34] , \sums[5][33] , \sums[5][32] , \sums[5][31] , \sums[5][30] , 
    \sums[5][29] , \sums[5][28] , \sums[5][27] , \sums[5][26] , \sums[5][25] , \sums[5][24] , 
    \sums[5][23] , \sums[5][22] , \sums[5][21] , \sums[5][20] , \sums[5][19] , \sums[5][18] , 
    \sums[5][17] , \sums[5][16] , uc_1286, uc_1287, uc_1288, uc_1289, uc_1290, uc_1291, 
    uc_1292, uc_1293, uc_1294, uc_1295, uc_1296, uc_1297, uc_1298, uc_1299, uc_1300, 
    uc_1301}), .v ({\couts[5][63] , uc_1302, uc_1303, uc_1304, uc_1305, uc_1306, 
    uc_1307, uc_1308, uc_1309, uc_1310, uc_1311, uc_1312, uc_1313, uc_1314, uc_1315, 
    \couts[5][48] , \couts[5][47] , \couts[5][46] , \couts[5][45] , \couts[5][44] , 
    \couts[5][43] , \couts[5][42] , \couts[5][41] , \couts[5][40] , \couts[5][39] , 
    \couts[5][38] , \couts[5][37] , \couts[5][36] , \couts[5][35] , \couts[5][34] , 
    \couts[5][33] , \couts[5][32] , \couts[5][31] , \couts[5][30] , \couts[5][29] , 
    \couts[5][28] , \couts[5][27] , \couts[5][26] , \couts[5][25] , \couts[5][24] , 
    \couts[5][23] , \couts[5][22] , \couts[5][21] , \couts[5][20] , \couts[5][19] , 
    \couts[5][18] , \couts[5][17] , uc_1316, uc_1317, uc_1318, uc_1319, uc_1320, 
    uc_1321, uc_1322, uc_1323, uc_1324, uc_1325, uc_1326, uc_1327, uc_1328, uc_1329, 
    uc_1330, uc_1331, uc_1332}), .x ({uc_1174, \pp[15][62] , uc_1175, uc_1176, uc_1177, 
    uc_1178, uc_1179, uc_1180, uc_1181, uc_1182, uc_1183, uc_1184, uc_1185, uc_1186, 
    uc_1187, uc_1188, uc_1189, uc_1190, \pp[15][45] , \pp[15][44] , \pp[15][43] , 
    \pp[15][42] , \pp[15][41] , \pp[15][40] , \pp[15][39] , \pp[15][38] , \pp[15][37] , 
    \pp[15][36] , \pp[15][35] , \pp[15][34] , \pp[15][33] , \pp[15][32] , \pp[15][31] , 
    \pp[15][30] , \pp[15][29] , \pp[15][28] , \pp[15][27] , \pp[15][26] , \pp[15][25] , 
    \pp[15][24] , \pp[15][23] , \pp[15][22] , \pp[15][21] , \pp[15][20] , \pp[15][19] , 
    \pp[15][18] , \pp[15][17] , \pp[15][16] , uc_1191, uc_1192, uc_1193, uc_1194, 
    uc_1195, uc_1196, uc_1197, uc_1198, uc_1199, uc_1200, uc_1201, uc_1202, uc_1203, 
    uc_1204, uc_1205, uc_1206}), .y ({uc_1207, \pp[16][62] , uc_1208, uc_1209, uc_1210, 
    uc_1211, uc_1212, uc_1213, uc_1214, uc_1215, uc_1216, uc_1217, uc_1218, uc_1219, 
    uc_1220, uc_1221, uc_1222, \pp[16][46] , \pp[16][45] , \pp[16][44] , \pp[16][43] , 
    \pp[16][42] , \pp[16][41] , \pp[16][40] , \pp[16][39] , \pp[16][38] , \pp[16][37] , 
    \pp[16][36] , \pp[16][35] , \pp[16][34] , \pp[16][33] , \pp[16][32] , \pp[16][31] , 
    \pp[16][30] , \pp[16][29] , \pp[16][28] , \pp[16][27] , \pp[16][26] , \pp[16][25] , 
    \pp[16][24] , \pp[16][23] , \pp[16][22] , \pp[16][21] , \pp[16][20] , \pp[16][19] , 
    \pp[16][18] , \pp[16][17] , \pp[16][16] , uc_1223, uc_1224, uc_1225, uc_1226, 
    uc_1227, uc_1228, uc_1229, uc_1230, uc_1231, uc_1232, uc_1233, uc_1234, uc_1235, 
    uc_1236, uc_1237, uc_1238}), .z ({uc_1239, \pp[17][62] , uc_1240, uc_1241, uc_1242, 
    uc_1243, uc_1244, uc_1245, uc_1246, uc_1247, uc_1248, uc_1249, uc_1250, uc_1251, 
    uc_1252, uc_1253, \pp[17][47] , \pp[17][46] , \pp[17][45] , \pp[17][44] , \pp[17][43] , 
    \pp[17][42] , \pp[17][41] , \pp[17][40] , \pp[17][39] , \pp[17][38] , \pp[17][37] , 
    \pp[17][36] , \pp[17][35] , \pp[17][34] , \pp[17][33] , \pp[17][32] , \pp[17][31] , 
    \pp[17][30] , \pp[17][29] , \pp[17][28] , \pp[17][27] , \pp[17][26] , \pp[17][25] , 
    \pp[17][24] , \pp[17][23] , \pp[17][22] , \pp[17][21] , \pp[17][20] , \pp[17][19] , 
    \pp[17][18] , \pp[17][17] , uc_1254, uc_1255, uc_1256, uc_1257, uc_1258, uc_1259, 
    uc_1260, uc_1261, uc_1262, uc_1263, uc_1264, uc_1265, uc_1266, uc_1267, uc_1268, 
    uc_1269, uc_1270}));
CSA__1_2 CSA13 (.u ({\sums[13][63] , uc_1116, uc_1117, uc_1118, uc_1119, uc_1120, 
    uc_1121, uc_1122, uc_1123, uc_1124, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, 
    \sums[13][48] , \sums[13][47] , \sums[13][46] , \sums[13][45] , \sums[13][44] , 
    \sums[13][43] , \sums[13][42] , \sums[13][41] , \sums[13][40] , \sums[13][39] , 
    \sums[13][38] , \sums[13][37] , \sums[13][36] , \sums[13][35] , \sums[13][34] , 
    \sums[13][33] , \sums[13][32] , \sums[13][31] , \sums[13][30] , \sums[13][29] , 
    \sums[13][28] , \sums[13][27] , \sums[13][26] , \sums[13][25] , \sums[13][24] , 
    \sums[13][23] , \sums[13][22] , \sums[13][21] , \sums[13][20] , \sums[13][19] , 
    \sums[13][18] , \sums[13][17] , \sums[13][16] , \sums[13][15] , uc_1130, uc_1131, 
    uc_1132, uc_1133, uc_1134, uc_1135, uc_1136, uc_1137, uc_1138, uc_1139, uc_1140, 
    uc_1141, uc_1142, uc_1143, uc_1144}), .v ({\couts[13][63] , uc_1145, uc_1146, 
    uc_1147, uc_1148, uc_1149, uc_1150, uc_1151, uc_1152, uc_1153, uc_1154, uc_1155, 
    uc_1156, uc_1157, \couts[13][49] , \couts[13][48] , \couts[13][47] , \couts[13][46] , 
    \couts[13][45] , \couts[13][44] , \couts[13][43] , \couts[13][42] , \couts[13][41] , 
    \couts[13][40] , \couts[13][39] , \couts[13][38] , \couts[13][37] , \couts[13][36] , 
    \couts[13][35] , \couts[13][34] , \couts[13][33] , \couts[13][32] , \couts[13][31] , 
    \couts[13][30] , \couts[13][29] , \couts[13][28] , \couts[13][27] , \couts[13][26] , 
    \couts[13][25] , \couts[13][24] , \couts[13][23] , \couts[13][22] , \couts[13][21] , 
    \couts[13][20] , \couts[13][19] , \couts[13][18] , \couts[13][17] , \couts[13][16] , 
    uc_1158, uc_1159, uc_1160, uc_1161, uc_1162, uc_1163, uc_1164, uc_1165, uc_1166, 
    uc_1167, uc_1168, uc_1169, uc_1170, uc_1171, uc_1172, uc_1173}), .x ({\couts[4][63] , 
    uc_1024, uc_1025, uc_1026, uc_1027, uc_1028, uc_1029, uc_1030, uc_1031, uc_1032, 
    uc_1033, uc_1034, uc_1035, uc_1036, uc_1037, uc_1038, uc_1039, uc_1040, \couts[4][45] , 
    \couts[4][44] , \couts[4][43] , \couts[4][42] , \couts[4][41] , \couts[4][40] , 
    \couts[4][39] , \couts[4][38] , \couts[4][37] , \couts[4][36] , \couts[4][35] , 
    \couts[4][34] , \couts[4][33] , \couts[4][32] , \couts[4][31] , \couts[4][30] , 
    \couts[4][29] , \couts[4][28] , \couts[4][27] , \couts[4][26] , \couts[4][25] , 
    \couts[4][24] , \couts[4][23] , \couts[4][22] , \couts[4][21] , \couts[4][20] , 
    \couts[4][19] , \couts[4][18] , \couts[4][17] , \couts[4][16] , \couts[4][15] , 
    uc_1041, uc_1042, uc_1043, uc_1044, uc_1045, uc_1046, uc_1047, uc_1048, uc_1049, 
    uc_1050, uc_1051, uc_1052, uc_1053, uc_1054, uc_1055}), .y ({\sums[5][63] , uc_1056, 
    uc_1057, uc_1058, uc_1059, uc_1060, uc_1061, uc_1062, uc_1063, uc_1064, uc_1065, 
    uc_1066, uc_1067, uc_1068, uc_1069, uc_1070, \sums[5][47] , \sums[5][46] , \sums[5][45] , 
    \sums[5][44] , \sums[5][43] , \sums[5][42] , \sums[5][41] , \sums[5][40] , \sums[5][39] , 
    \sums[5][38] , \sums[5][37] , \sums[5][36] , \sums[5][35] , \sums[5][34] , \sums[5][33] , 
    \sums[5][32] , \sums[5][31] , \sums[5][30] , \sums[5][29] , \sums[5][28] , \sums[5][27] , 
    \sums[5][26] , \sums[5][25] , \sums[5][24] , \sums[5][23] , \sums[5][22] , \sums[5][21] , 
    \sums[5][20] , \sums[5][19] , \sums[5][18] , \sums[5][17] , \sums[5][16] , \pp[15][15] , 
    uc_1071, uc_1072, uc_1073, uc_1074, uc_1075, uc_1076, uc_1077, uc_1078, uc_1079, 
    uc_1080, uc_1081, uc_1082, uc_1083, uc_1084, 1'b0 }), .z ({\couts[5][63] , uc_1085, 
    uc_1086, uc_1087, uc_1088, uc_1089, uc_1090, uc_1091, uc_1092, uc_1093, uc_1094, 
    uc_1095, uc_1096, uc_1097, uc_1098, \couts[5][48] , \couts[5][47] , \couts[5][46] , 
    \couts[5][45] , \couts[5][44] , \couts[5][43] , \couts[5][42] , \couts[5][41] , 
    \couts[5][40] , \couts[5][39] , \couts[5][38] , \couts[5][37] , \couts[5][36] , 
    \couts[5][35] , \couts[5][34] , \couts[5][33] , \couts[5][32] , \couts[5][31] , 
    \couts[5][30] , \couts[5][29] , \couts[5][28] , \couts[5][27] , \couts[5][26] , 
    \couts[5][25] , \couts[5][24] , \couts[5][23] , \couts[5][22] , \couts[5][21] , 
    \couts[5][20] , \couts[5][19] , \couts[5][18] , \couts[5][17] , uc_1099, uc_1100, 
    uc_1101, uc_1102, uc_1103, uc_1104, uc_1105, uc_1106, uc_1107, uc_1108, uc_1109, 
    uc_1110, uc_1111, uc_1112, uc_1113, uc_1114, uc_1115}));
products Products (.\pp[0]  ({\pp[0][63] , uc_992, uc_993, uc_994, uc_995, uc_996, 
    uc_997, uc_998, uc_999, uc_1000, uc_1001, uc_1002, uc_1003, uc_1004, uc_1005, 
    uc_1006, uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, uc_1013, uc_1014, 
    uc_1015, uc_1016, uc_1017, uc_1018, uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, 
    \pp[0][30] , \pp[0][29] , \pp[0][28] , \pp[0][27] , \pp[0][26] , \pp[0][25] , 
    \pp[0][24] , \pp[0][23] , \pp[0][22] , \pp[0][21] , \pp[0][20] , \pp[0][19] , 
    \pp[0][18] , \pp[0][17] , \pp[0][16] , \pp[0][15] , \pp[0][14] , \pp[0][13] , 
    \pp[0][12] , \pp[0][11] , \pp[0][10] , \pp[0][9] , \pp[0][8] , \pp[0][7] , \pp[0][6] , 
    \pp[0][5] , \pp[0][4] , \pp[0][3] , \pp[0][2] , \pp[0][1] , out[0]}), .\pp[10]  ({
    \pp[10][63] , uc_672, uc_673, uc_674, uc_675, uc_676, uc_677, uc_678, uc_679, 
    uc_680, uc_681, uc_682, uc_683, uc_684, uc_685, uc_686, uc_687, uc_688, uc_689, 
    uc_690, uc_691, uc_692, uc_693, \pp[10][40] , \pp[10][39] , \pp[10][38] , \pp[10][37] , 
    \pp[10][36] , \pp[10][35] , \pp[10][34] , \pp[10][33] , \pp[10][32] , \pp[10][31] , 
    \pp[10][30] , \pp[10][29] , \pp[10][28] , \pp[10][27] , \pp[10][26] , \pp[10][25] , 
    \pp[10][24] , \pp[10][23] , \pp[10][22] , \pp[10][21] , \pp[10][20] , \pp[10][19] , 
    \pp[10][18] , \pp[10][17] , \pp[10][16] , \pp[10][15] , \pp[10][14] , \pp[10][13] , 
    \pp[10][12] , \pp[10][11] , \pp[10][10] , uc_694, uc_695, uc_696, uc_697, uc_698, 
    uc_699, uc_700, uc_701, uc_702, uc_703}), .\pp[11]  ({\pp[11][63] , uc_640, uc_641, 
    uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, uc_651, 
    uc_652, uc_653, uc_654, uc_655, uc_656, uc_657, uc_658, uc_659, uc_660, \pp[11][41] , 
    \pp[11][40] , \pp[11][39] , \pp[11][38] , \pp[11][37] , \pp[11][36] , \pp[11][35] , 
    \pp[11][34] , \pp[11][33] , \pp[11][32] , \pp[11][31] , \pp[11][30] , \pp[11][29] , 
    \pp[11][28] , \pp[11][27] , \pp[11][26] , \pp[11][25] , \pp[11][24] , \pp[11][23] , 
    \pp[11][22] , \pp[11][21] , \pp[11][20] , \pp[11][19] , \pp[11][18] , \pp[11][17] , 
    \pp[11][16] , \pp[11][15] , \pp[11][14] , \pp[11][13] , \pp[11][12] , \pp[11][11] , 
    uc_661, uc_662, uc_663, uc_664, uc_665, uc_666, uc_667, uc_668, uc_669, uc_670, 
    uc_671}), .\pp[12]  ({uc_608, \pp[12][62] , uc_609, uc_610, uc_611, uc_612, uc_613, 
    uc_614, uc_615, uc_616, uc_617, uc_618, uc_619, uc_620, uc_621, uc_622, uc_623, 
    uc_624, uc_625, uc_626, uc_627, \pp[12][42] , \pp[12][41] , \pp[12][40] , \pp[12][39] , 
    \pp[12][38] , \pp[12][37] , \pp[12][36] , \pp[12][35] , \pp[12][34] , \pp[12][33] , 
    \pp[12][32] , \pp[12][31] , \pp[12][30] , \pp[12][29] , \pp[12][28] , \pp[12][27] , 
    \pp[12][26] , \pp[12][25] , \pp[12][24] , \pp[12][23] , \pp[12][22] , \pp[12][21] , 
    \pp[12][20] , \pp[12][19] , \pp[12][18] , \pp[12][17] , \pp[12][16] , \pp[12][15] , 
    \pp[12][14] , \pp[12][13] , \sums[4][12] , uc_628, uc_629, uc_630, uc_631, uc_632, 
    uc_633, uc_634, uc_635, uc_636, uc_637, uc_638, uc_639}), .\pp[13]  ({uc_576, 
    \pp[13][62] , uc_577, uc_578, uc_579, uc_580, uc_581, uc_582, uc_583, uc_584, 
    uc_585, uc_586, uc_587, uc_588, uc_589, uc_590, uc_591, uc_592, uc_593, uc_594, 
    \pp[13][43] , \pp[13][42] , \pp[13][41] , \pp[13][40] , \pp[13][39] , \pp[13][38] , 
    \pp[13][37] , \pp[13][36] , \pp[13][35] , \pp[13][34] , \pp[13][33] , \pp[13][32] , 
    \pp[13][31] , \pp[13][30] , \pp[13][29] , \pp[13][28] , \pp[13][27] , \pp[13][26] , 
    \pp[13][25] , \pp[13][24] , \pp[13][23] , \pp[13][22] , \pp[13][21] , \pp[13][20] , 
    \pp[13][19] , \pp[13][18] , \pp[13][17] , \pp[13][16] , \pp[13][15] , \pp[13][14] , 
    \pp[13][13] , uc_595, uc_596, uc_597, uc_598, uc_599, uc_600, uc_601, uc_602, 
    uc_603, uc_604, uc_605, uc_606, uc_607}), .\pp[14]  ({uc_544, \pp[14][62] , uc_545, 
    uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, uc_555, 
    uc_556, uc_557, uc_558, uc_559, uc_560, uc_561, \pp[14][44] , \pp[14][43] , \pp[14][42] , 
    \pp[14][41] , \pp[14][40] , \pp[14][39] , \pp[14][38] , \pp[14][37] , \pp[14][36] , 
    \pp[14][35] , \pp[14][34] , \pp[14][33] , \pp[14][32] , \pp[14][31] , \pp[14][30] , 
    \pp[14][29] , \pp[14][28] , \pp[14][27] , \pp[14][26] , \pp[14][25] , \pp[14][24] , 
    \pp[14][23] , \pp[14][22] , \pp[14][21] , \pp[14][20] , \pp[14][19] , \pp[14][18] , 
    \pp[14][17] , \pp[14][16] , \pp[14][15] , \pp[14][14] , uc_562, uc_563, uc_564, 
    uc_565, uc_566, uc_567, uc_568, uc_569, uc_570, uc_571, uc_572, uc_573, uc_574, 
    uc_575}), .\pp[15]  ({uc_512, \pp[15][62] , uc_513, uc_514, uc_515, uc_516, uc_517, 
    uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, uc_525, uc_526, uc_527, 
    uc_528, \pp[15][45] , \pp[15][44] , \pp[15][43] , \pp[15][42] , \pp[15][41] , 
    \pp[15][40] , \pp[15][39] , \pp[15][38] , \pp[15][37] , \pp[15][36] , \pp[15][35] , 
    \pp[15][34] , \pp[15][33] , \pp[15][32] , \pp[15][31] , \pp[15][30] , \pp[15][29] , 
    \pp[15][28] , \pp[15][27] , \pp[15][26] , \pp[15][25] , \pp[15][24] , \pp[15][23] , 
    \pp[15][22] , \pp[15][21] , \pp[15][20] , \pp[15][19] , \pp[15][18] , \pp[15][17] , 
    \pp[15][16] , \pp[15][15] , uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, uc_535, 
    uc_536, uc_537, uc_538, uc_539, uc_540, uc_541, uc_542, uc_543}), .\pp[16]  ({
    uc_480, \pp[16][62] , uc_481, uc_482, uc_483, uc_484, uc_485, uc_486, uc_487, 
    uc_488, uc_489, uc_490, uc_491, uc_492, uc_493, uc_494, uc_495, \pp[16][46] , 
    \pp[16][45] , \pp[16][44] , \pp[16][43] , \pp[16][42] , \pp[16][41] , \pp[16][40] , 
    \pp[16][39] , \pp[16][38] , \pp[16][37] , \pp[16][36] , \pp[16][35] , \pp[16][34] , 
    \pp[16][33] , \pp[16][32] , \pp[16][31] , \pp[16][30] , \pp[16][29] , \pp[16][28] , 
    \pp[16][27] , \pp[16][26] , \pp[16][25] , \pp[16][24] , \pp[16][23] , \pp[16][22] , 
    \pp[16][21] , \pp[16][20] , \pp[16][19] , \pp[16][18] , \pp[16][17] , \pp[16][16] , 
    uc_496, uc_497, uc_498, uc_499, uc_500, uc_501, uc_502, uc_503, uc_504, uc_505, 
    uc_506, uc_507, uc_508, uc_509, uc_510, uc_511}), .\pp[17]  ({uc_448, \pp[17][62] , 
    uc_449, uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, 
    uc_459, uc_460, uc_461, uc_462, \pp[17][47] , \pp[17][46] , \pp[17][45] , \pp[17][44] , 
    \pp[17][43] , \pp[17][42] , \pp[17][41] , \pp[17][40] , \pp[17][39] , \pp[17][38] , 
    \pp[17][37] , \pp[17][36] , \pp[17][35] , \pp[17][34] , \pp[17][33] , \pp[17][32] , 
    \pp[17][31] , \pp[17][30] , \pp[17][29] , \pp[17][28] , \pp[17][27] , \pp[17][26] , 
    \pp[17][25] , \pp[17][24] , \pp[17][23] , \pp[17][22] , \pp[17][21] , \pp[17][20] , 
    \pp[17][19] , \pp[17][18] , \pp[17][17] , uc_463, uc_464, uc_465, uc_466, uc_467, 
    uc_468, uc_469, uc_470, uc_471, uc_472, uc_473, uc_474, uc_475, uc_476, uc_477, 
    uc_478, uc_479}), .\pp[18]  ({\pp[18][63] , uc_416, uc_417, uc_418, uc_419, uc_420, 
    uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, uc_429, \pp[18][48] , 
    \pp[18][47] , \pp[18][46] , \pp[18][45] , \pp[18][44] , \pp[18][43] , \pp[18][42] , 
    \pp[18][41] , \pp[18][40] , \pp[18][39] , \pp[18][38] , \pp[18][37] , \pp[18][36] , 
    \pp[18][35] , \pp[18][34] , \pp[18][33] , \pp[18][32] , \pp[18][31] , \pp[18][30] , 
    \pp[18][29] , \pp[18][28] , \pp[18][27] , \pp[18][26] , \pp[18][25] , \pp[18][24] , 
    \pp[18][23] , \pp[18][22] , \pp[18][21] , \pp[18][20] , \pp[18][19] , \pp[18][18] , 
    uc_430, uc_431, uc_432, uc_433, uc_434, uc_435, uc_436, uc_437, uc_438, uc_439, 
    uc_440, uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, uc_447}), .\pp[19]  ({
    \pp[19][63] , uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, uc_390, uc_391, 
    uc_392, uc_393, uc_394, uc_395, uc_396, \pp[19][49] , \pp[19][48] , \pp[19][47] , 
    \pp[19][46] , \pp[19][45] , \pp[19][44] , \pp[19][43] , \pp[19][42] , \pp[19][41] , 
    \pp[19][40] , \pp[19][39] , \pp[19][38] , \pp[19][37] , \pp[19][36] , \pp[19][35] , 
    \pp[19][34] , \pp[19][33] , \pp[19][32] , \pp[19][31] , \pp[19][30] , \pp[19][29] , 
    \pp[19][28] , \pp[19][27] , \pp[19][26] , \pp[19][25] , \pp[19][24] , \pp[19][23] , 
    \pp[19][22] , \pp[19][21] , \pp[19][20] , \pp[19][19] , uc_397, uc_398, uc_399, 
    uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, uc_408, uc_409, 
    uc_410, uc_411, uc_412, uc_413, uc_414, uc_415}), .\pp[1]  ({\pp[1][63] , uc_960, 
    uc_961, uc_962, uc_963, uc_964, uc_965, uc_966, uc_967, uc_968, uc_969, uc_970, 
    uc_971, uc_972, uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, uc_979, uc_980, 
    uc_981, uc_982, uc_983, uc_984, uc_985, uc_986, uc_987, uc_988, uc_989, uc_990, 
    \pp[1][31] , \pp[1][30] , \pp[1][29] , \pp[1][28] , \pp[1][27] , \pp[1][26] , 
    \pp[1][25] , \pp[1][24] , \pp[1][23] , \pp[1][22] , \pp[1][21] , \pp[1][20] , 
    \pp[1][19] , \pp[1][18] , \pp[1][17] , \pp[1][16] , \pp[1][15] , \pp[1][14] , 
    \pp[1][13] , \pp[1][12] , \pp[1][11] , \pp[1][10] , \pp[1][9] , \pp[1][8] , \pp[1][7] , 
    \pp[1][6] , \pp[1][5] , \pp[1][4] , \pp[1][3] , \pp[1][2] , \pp[1][1] , uc_991})
    , .\pp[20]  ({\pp[20][63] , uc_352, uc_353, uc_354, uc_355, uc_356, uc_357, uc_358, 
    uc_359, uc_360, uc_361, uc_362, uc_363, \pp[20][50] , \pp[20][49] , \pp[20][48] , 
    \pp[20][47] , \pp[20][46] , \pp[20][45] , \pp[20][44] , \pp[20][43] , \pp[20][42] , 
    \pp[20][41] , \pp[20][40] , \pp[20][39] , \pp[20][38] , \pp[20][37] , \pp[20][36] , 
    \pp[20][35] , \pp[20][34] , \pp[20][33] , \pp[20][32] , \pp[20][31] , \pp[20][30] , 
    \pp[20][29] , \pp[20][28] , \pp[20][27] , \pp[20][26] , \pp[20][25] , \pp[20][24] , 
    \pp[20][23] , \pp[20][22] , \pp[20][21] , \pp[20][20] , uc_364, uc_365, uc_366, 
    uc_367, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374, uc_375, uc_376, 
    uc_377, uc_378, uc_379, uc_380, uc_381, uc_382, uc_383}), .\pp[21]  ({\pp[21][63] , 
    uc_320, uc_321, uc_322, uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, 
    uc_330, \pp[21][51] , \pp[21][50] , \pp[21][49] , \pp[21][48] , \pp[21][47] , 
    \pp[21][46] , \pp[21][45] , \pp[21][44] , \pp[21][43] , \pp[21][42] , \pp[21][41] , 
    \pp[21][40] , \pp[21][39] , \pp[21][38] , \pp[21][37] , \pp[21][36] , \pp[21][35] , 
    \pp[21][34] , \pp[21][33] , \pp[21][32] , \pp[21][31] , \pp[21][30] , \pp[21][29] , 
    \pp[21][28] , \pp[21][27] , \pp[21][26] , \pp[21][25] , \pp[21][24] , \pp[21][23] , 
    \pp[21][22] , \pp[21][21] , uc_331, uc_332, uc_333, uc_334, uc_335, uc_336, uc_337, 
    uc_338, uc_339, uc_340, uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, 
    uc_348, uc_349, uc_350, uc_351}), .\pp[22]  ({\pp[22][63] , uc_288, uc_289, uc_290, 
    uc_291, uc_292, uc_293, uc_294, uc_295, uc_296, uc_297, \pp[22][52] , \pp[22][51] , 
    \pp[22][50] , \pp[22][49] , \pp[22][48] , \pp[22][47] , \pp[22][46] , \pp[22][45] , 
    \pp[22][44] , \pp[22][43] , \pp[22][42] , \pp[22][41] , \pp[22][40] , \pp[22][39] , 
    \pp[22][38] , \pp[22][37] , \pp[22][36] , \pp[22][35] , \pp[22][34] , \pp[22][33] , 
    \pp[22][32] , \pp[22][31] , \pp[22][30] , \pp[22][29] , \pp[22][28] , \pp[22][27] , 
    \pp[22][26] , \pp[22][25] , \pp[22][24] , \pp[22][23] , \pp[22][22] , uc_298, 
    uc_299, uc_300, uc_301, uc_302, uc_303, uc_304, uc_305, uc_306, uc_307, uc_308, 
    uc_309, uc_310, uc_311, uc_312, uc_313, uc_314, uc_315, uc_316, uc_317, uc_318, 
    uc_319}), .\pp[23]  ({\pp[23][63] , uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, 
    uc_262, uc_263, uc_264, \pp[23][53] , \pp[23][52] , \pp[23][51] , \pp[23][50] , 
    \pp[23][49] , \pp[23][48] , \pp[23][47] , \pp[23][46] , \pp[23][45] , \pp[23][44] , 
    \pp[23][43] , \pp[23][42] , \pp[23][41] , \pp[23][40] , \pp[23][39] , \pp[23][38] , 
    \pp[23][37] , \pp[23][36] , \pp[23][35] , \pp[23][34] , \pp[23][33] , \pp[23][32] , 
    \pp[23][31] , \pp[23][30] , \pp[23][29] , \pp[23][28] , \pp[23][27] , \pp[23][26] , 
    \pp[23][25] , \pp[23][24] , \pp[23][23] , uc_265, uc_266, uc_267, uc_268, uc_269, 
    uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, uc_276, uc_277, uc_278, uc_279, 
    uc_280, uc_281, uc_282, uc_283, uc_284, uc_285, uc_286, uc_287}), .\pp[24]  ({
    \pp[24][63] , uc_224, uc_225, uc_226, uc_227, uc_228, uc_229, uc_230, uc_231, 
    \pp[24][54] , \pp[24][53] , \pp[24][52] , \pp[24][51] , \pp[24][50] , \pp[24][49] , 
    \pp[24][48] , \pp[24][47] , \pp[24][46] , \pp[24][45] , \pp[24][44] , \pp[24][43] , 
    \pp[24][42] , \pp[24][41] , \pp[24][40] , \pp[24][39] , \pp[24][38] , \pp[24][37] , 
    \pp[24][36] , \pp[24][35] , \pp[24][34] , \pp[24][33] , \pp[24][32] , \pp[24][31] , 
    \pp[24][30] , \pp[24][29] , \pp[24][28] , \pp[24][27] , \pp[24][26] , \pp[24][25] , 
    \pp[24][24] , uc_232, uc_233, uc_234, uc_235, uc_236, uc_237, uc_238, uc_239, 
    uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, uc_247, uc_248, uc_249, 
    uc_250, uc_251, uc_252, uc_253, uc_254, uc_255}), .\pp[25]  ({\pp[25][63] , uc_192, 
    uc_193, uc_194, uc_195, uc_196, uc_197, uc_198, \pp[25][55] , \pp[25][54] , \pp[25][53] , 
    \pp[25][52] , \pp[25][51] , \pp[25][50] , \pp[25][49] , \pp[25][48] , \pp[25][47] , 
    \pp[25][46] , \pp[25][45] , \pp[25][44] , \pp[25][43] , \pp[25][42] , \pp[25][41] , 
    \pp[25][40] , \pp[25][39] , \pp[25][38] , \pp[25][37] , \pp[25][36] , \pp[25][35] , 
    \pp[25][34] , \pp[25][33] , \pp[25][32] , \pp[25][31] , \pp[25][30] , \pp[25][29] , 
    \pp[25][28] , \pp[25][27] , \pp[25][26] , \pp[25][25] , uc_199, uc_200, uc_201, 
    uc_202, uc_203, uc_204, uc_205, uc_206, uc_207, uc_208, uc_209, uc_210, uc_211, 
    uc_212, uc_213, uc_214, uc_215, uc_216, uc_217, uc_218, uc_219, uc_220, uc_221, 
    uc_222, uc_223}), .\pp[26]  ({\pp[26][63] , uc_160, uc_161, uc_162, uc_163, uc_164, 
    uc_165, \pp[26][56] , \pp[26][55] , \pp[26][54] , \pp[26][53] , \pp[26][52] , 
    \pp[26][51] , \pp[26][50] , \pp[26][49] , \pp[26][48] , \pp[26][47] , \pp[26][46] , 
    \pp[26][45] , \pp[26][44] , \pp[26][43] , \pp[26][42] , \pp[26][41] , \pp[26][40] , 
    \pp[26][39] , \pp[26][38] , \pp[26][37] , \pp[26][36] , \pp[26][35] , \pp[26][34] , 
    \pp[26][33] , \pp[26][32] , \pp[26][31] , \pp[26][30] , \pp[26][29] , \pp[26][28] , 
    \pp[26][27] , \pp[26][26] , uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, uc_172, 
    uc_173, uc_174, uc_175, uc_176, uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, 
    uc_183, uc_184, uc_185, uc_186, uc_187, uc_188, uc_189, uc_190, uc_191}), .\pp[27]  ({
    \pp[27][58] , uc_128, uc_129, uc_130, uc_131, uc_132, \pp[27][57] , \pp[27][56] , 
    \pp[27][55] , \pp[27][54] , \pp[27][53] , \pp[27][52] , \pp[27][51] , \pp[27][50] , 
    \pp[27][49] , \pp[27][48] , \pp[27][47] , \pp[27][46] , \pp[27][45] , \pp[27][44] , 
    \pp[27][43] , \pp[27][42] , \pp[27][41] , \pp[27][40] , \pp[27][39] , \pp[27][38] , 
    \pp[27][37] , \pp[27][36] , \pp[27][35] , \pp[27][34] , \pp[27][33] , \pp[27][32] , 
    \pp[27][31] , \pp[27][30] , \pp[27][29] , \pp[27][28] , \pp[27][27] , uc_133, 
    uc_134, uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, 
    uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, uc_153, 
    uc_154, uc_155, uc_156, uc_157, uc_158, uc_159}), .\pp[28]  ({\pp[28][63] , uc_96, 
    uc_97, uc_98, uc_99, \pp[28][58] , \pp[28][57] , \pp[28][56] , \pp[28][55] , 
    \pp[28][54] , \pp[28][53] , \pp[28][52] , \pp[28][51] , \pp[28][50] , \pp[28][49] , 
    \pp[28][48] , \pp[28][47] , \pp[28][46] , \pp[28][45] , \pp[28][44] , \pp[28][43] , 
    \pp[28][42] , \pp[28][41] , \pp[28][40] , \pp[28][39] , \pp[28][38] , \pp[28][37] , 
    \pp[28][36] , \pp[28][35] , \pp[28][34] , \pp[28][33] , \pp[28][32] , \pp[28][31] , 
    \pp[28][30] , \pp[28][29] , \pp[28][28] , uc_100, uc_101, uc_102, uc_103, uc_104, 
    uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, 
    uc_115, uc_116, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, uc_124, 
    uc_125, uc_126, uc_127}), .\pp[29]  ({\pp[29][63] , uc_64, uc_65, uc_66, \pp[29][59] , 
    \pp[29][58] , \pp[29][57] , \pp[29][56] , \pp[29][55] , \pp[29][54] , \pp[29][53] , 
    \pp[29][52] , \pp[29][51] , \pp[29][50] , \pp[29][49] , \pp[29][48] , \pp[29][47] , 
    \pp[29][46] , \pp[29][45] , \pp[29][44] , \pp[29][43] , \pp[29][42] , \pp[29][41] , 
    \pp[29][40] , \pp[29][39] , \pp[29][38] , \pp[29][37] , \pp[29][36] , \pp[29][35] , 
    \pp[29][34] , \pp[29][33] , \pp[29][32] , \pp[29][31] , \pp[29][30] , \pp[29][29] , 
    uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, 
    uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, 
    uc_89, uc_90, uc_91, uc_92, uc_93, uc_94, uc_95}), .\pp[2]  ({\pp[2][63] , uc_928, 
    uc_929, uc_930, uc_931, uc_932, uc_933, uc_934, uc_935, uc_936, uc_937, uc_938, 
    uc_939, uc_940, uc_941, uc_942, uc_943, uc_944, uc_945, uc_946, uc_947, uc_948, 
    uc_949, uc_950, uc_951, uc_952, uc_953, uc_954, uc_955, uc_956, uc_957, \pp[2][32] , 
    \pp[2][31] , \pp[2][30] , \pp[2][29] , \pp[2][28] , \pp[2][27] , \pp[2][26] , 
    \pp[2][25] , \pp[2][24] , \pp[2][23] , \pp[2][22] , \pp[2][21] , \pp[2][20] , 
    \pp[2][19] , \pp[2][18] , \pp[2][17] , \pp[2][16] , \pp[2][15] , \pp[2][14] , 
    \pp[2][13] , \pp[2][12] , \pp[2][11] , \pp[2][10] , \pp[2][9] , \pp[2][8] , \pp[2][7] , 
    \pp[2][6] , \pp[2][5] , \pp[2][4] , \pp[2][3] , \pp[2][2] , uc_958, uc_959}), .\pp[30]  ({
    \pp[30][63] , uc_32, uc_33, \pp[30][60] , \pp[30][59] , \pp[30][58] , \pp[30][57] , 
    \pp[30][56] , \pp[30][55] , \pp[30][54] , \pp[30][53] , \pp[30][52] , \pp[30][51] , 
    \pp[30][50] , \pp[30][49] , \pp[30][48] , \pp[30][47] , \pp[30][46] , \pp[30][45] , 
    \pp[30][44] , \pp[30][43] , \pp[30][42] , \pp[30][41] , \pp[30][40] , \pp[30][39] , 
    \pp[30][38] , \pp[30][37] , \pp[30][36] , \pp[30][35] , \pp[30][34] , \pp[30][33] , 
    \pp[30][32] , \pp[30][31] , \pp[30][30] , uc_34, uc_35, uc_36, uc_37, uc_38, 
    uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, 
    uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, 
    uc_61, uc_62, uc_63}), .\pp[31]  ({\pp[31][63] , uc_0, \pp[31][61] , \pp[31][60] , 
    \pp[31][59] , \pp[31][58] , \pp[31][57] , \pp[31][56] , \pp[31][55] , \pp[31][54] , 
    \pp[31][53] , \pp[31][52] , \pp[31][51] , \pp[31][50] , \pp[31][49] , \pp[31][48] , 
    \pp[31][47] , \pp[31][46] , \pp[31][45] , \pp[31][44] , \pp[31][43] , \pp[31][42] , 
    \pp[31][41] , \pp[31][40] , \pp[31][39] , \pp[31][38] , \pp[31][37] , \pp[31][36] , 
    \pp[31][35] , \pp[31][34] , \pp[31][33] , \pp[31][32] , \pp[31][31] , uc_1, uc_2, 
    uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, 
    uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, 
    uc_26, uc_27, uc_28, uc_29, uc_30, uc_31}), .\pp[3]  ({\pp[3][63] , uc_896, uc_897, 
    uc_898, uc_899, uc_900, uc_901, uc_902, uc_903, uc_904, uc_905, uc_906, uc_907, 
    uc_908, uc_909, uc_910, uc_911, uc_912, uc_913, uc_914, uc_915, uc_916, uc_917, 
    uc_918, uc_919, uc_920, uc_921, uc_922, uc_923, uc_924, \pp[3][33] , \pp[3][32] , 
    \pp[3][31] , \pp[3][30] , \pp[3][29] , \pp[3][28] , \pp[3][27] , \pp[3][26] , 
    \pp[3][25] , \pp[3][24] , \pp[3][23] , \pp[3][22] , \pp[3][21] , \pp[3][20] , 
    \pp[3][19] , \pp[3][18] , \pp[3][17] , \pp[3][16] , \pp[3][15] , \pp[3][14] , 
    \pp[3][13] , \pp[3][12] , \pp[3][11] , \pp[3][10] , \pp[3][9] , \pp[3][8] , \pp[3][7] , 
    \pp[3][6] , \pp[3][5] , \pp[3][4] , \pp[3][3] , uc_925, uc_926, uc_927}), .\pp[4]  ({
    \pp[4][63] , uc_864, uc_865, uc_866, uc_867, uc_868, uc_869, uc_870, uc_871, 
    uc_872, uc_873, uc_874, uc_875, uc_876, uc_877, uc_878, uc_879, uc_880, uc_881, 
    uc_882, uc_883, uc_884, uc_885, uc_886, uc_887, uc_888, uc_889, uc_890, uc_891, 
    \pp[4][34] , \pp[4][33] , \pp[4][32] , \pp[4][31] , \pp[4][30] , \pp[4][29] , 
    \pp[4][28] , \pp[4][27] , \pp[4][26] , \pp[4][25] , \pp[4][24] , \pp[4][23] , 
    \pp[4][22] , \pp[4][21] , \pp[4][20] , \pp[4][19] , \pp[4][18] , \pp[4][17] , 
    \pp[4][16] , \pp[4][15] , \pp[4][14] , \pp[4][13] , \pp[4][12] , \pp[4][11] , 
    \pp[4][10] , \pp[4][9] , \pp[4][8] , \pp[4][7] , \pp[4][6] , \pp[4][5] , \pp[4][4] , 
    uc_892, uc_893, uc_894, uc_895}), .\pp[5]  ({\pp[5][63] , uc_832, uc_833, uc_834, 
    uc_835, uc_836, uc_837, uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, uc_844, 
    uc_845, uc_846, uc_847, uc_848, uc_849, uc_850, uc_851, uc_852, uc_853, uc_854, 
    uc_855, uc_856, uc_857, uc_858, \pp[5][35] , \pp[5][34] , \pp[5][33] , \pp[5][32] , 
    \pp[5][31] , \pp[5][30] , \pp[5][29] , \pp[5][28] , \pp[5][27] , \pp[5][26] , 
    \pp[5][25] , \pp[5][24] , \pp[5][23] , \pp[5][22] , \pp[5][21] , \pp[5][20] , 
    \pp[5][19] , \pp[5][18] , \pp[5][17] , \pp[5][16] , \pp[5][15] , \pp[5][14] , 
    \pp[5][13] , \pp[5][12] , \pp[5][11] , \pp[5][10] , \pp[5][9] , \pp[5][8] , \pp[5][7] , 
    \pp[5][6] , \pp[5][5] , uc_859, uc_860, uc_861, uc_862, uc_863}), .\pp[6]  ({
    \pp[6][63] , uc_800, uc_801, uc_802, uc_803, uc_804, uc_805, uc_806, uc_807, 
    uc_808, uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, uc_816, uc_817, 
    uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, \pp[6][36] , 
    \pp[6][35] , \pp[6][34] , \pp[6][33] , \pp[6][32] , \pp[6][31] , \pp[6][30] , 
    \pp[6][29] , \pp[6][28] , \pp[6][27] , \pp[6][26] , \pp[6][25] , \pp[6][24] , 
    \pp[6][23] , \pp[6][22] , \pp[6][21] , \pp[6][20] , \pp[6][19] , \pp[6][18] , 
    \pp[6][17] , \pp[6][16] , \pp[6][15] , \pp[6][14] , \pp[6][13] , \pp[6][12] , 
    \pp[6][11] , \pp[6][10] , \pp[6][9] , \pp[6][8] , \pp[6][7] , \pp[6][6] , uc_826, 
    uc_827, uc_828, uc_829, uc_830, uc_831}), .\pp[7]  ({\pp[7][63] , uc_768, uc_769, 
    uc_770, uc_771, uc_772, uc_773, uc_774, uc_775, uc_776, uc_777, uc_778, uc_779, 
    uc_780, uc_781, uc_782, uc_783, uc_784, uc_785, uc_786, uc_787, uc_788, uc_789, 
    uc_790, uc_791, uc_792, \pp[7][37] , \pp[7][36] , \pp[7][35] , \pp[7][34] , \pp[7][33] , 
    \pp[7][32] , \pp[7][31] , \pp[7][30] , \pp[7][29] , \pp[7][28] , \pp[7][27] , 
    \pp[7][26] , \pp[7][25] , \pp[7][24] , \pp[7][23] , \pp[7][22] , \pp[7][21] , 
    \pp[7][20] , \pp[7][19] , \pp[7][18] , \pp[7][17] , \pp[7][16] , \pp[7][15] , 
    \pp[7][14] , \pp[7][13] , \pp[7][12] , \pp[7][11] , \pp[7][10] , \pp[7][9] , 
    \pp[7][8] , \pp[7][7] , uc_793, uc_794, uc_795, uc_796, uc_797, uc_798, uc_799})
    , .\pp[8]  ({\pp[8][63] , uc_736, uc_737, uc_738, uc_739, uc_740, uc_741, uc_742, 
    uc_743, uc_744, uc_745, uc_746, uc_747, uc_748, uc_749, uc_750, uc_751, uc_752, 
    uc_753, uc_754, uc_755, uc_756, uc_757, uc_758, uc_759, \pp[8][38] , \pp[8][37] , 
    \pp[8][36] , \pp[8][35] , \pp[8][34] , \pp[8][33] , \pp[8][32] , \pp[8][31] , 
    \pp[8][30] , \pp[8][29] , \pp[8][28] , \pp[8][27] , \pp[8][26] , \pp[8][25] , 
    \pp[8][24] , \pp[8][23] , \pp[8][22] , \pp[8][21] , \pp[8][20] , \pp[8][19] , 
    \pp[8][18] , \pp[8][17] , \pp[8][16] , \pp[8][15] , \pp[8][14] , \pp[8][13] , 
    \pp[8][12] , \pp[8][11] , \pp[8][10] , \pp[8][9] , \pp[8][8] , uc_760, uc_761, 
    uc_762, uc_763, uc_764, uc_765, uc_766, uc_767}), .\pp[9]  ({\pp[9][63] , uc_704, 
    uc_705, uc_706, uc_707, uc_708, uc_709, uc_710, uc_711, uc_712, uc_713, uc_714, 
    uc_715, uc_716, uc_717, uc_718, uc_719, uc_720, uc_721, uc_722, uc_723, uc_724, 
    uc_725, uc_726, \pp[9][39] , \pp[9][38] , \pp[9][37] , \pp[9][36] , \pp[9][35] , 
    \pp[9][34] , \pp[9][33] , \pp[9][32] , \pp[9][31] , \pp[9][30] , \pp[9][29] , 
    \pp[9][28] , \pp[9][27] , \pp[9][26] , \pp[9][25] , \pp[9][24] , \pp[9][23] , 
    \pp[9][22] , \pp[9][21] , \pp[9][20] , \pp[9][19] , \pp[9][18] , \pp[9][17] , 
    \pp[9][16] , \pp[9][15] , \pp[9][14] , \pp[9][13] , \pp[9][12] , \pp[9][11] , 
    \pp[9][10] , \pp[9][9] , uc_727, uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, 
    uc_734, uc_735}), .x ({x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], 
    x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], 
    x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]})
    , .y ({y[31], y[30], y[29], y[28], y[27], y[26], y[25], y[24], y[23], y[22], 
    y[21], y[20], y[19], y[18], y[17], y[16], y[15], y[14], y[13], y[12], y[11], 
    y[10], y[9], y[8], y[7], y[6], y[5], y[4], y[3], y[2], y[1], y[0]}));

endmodule //mulTree

module integrationMult (clk, reset, en, inputA, inputB, result);

output [63:0] result;
input clk;
input en;
input [31:0] inputA;
input [31:0] inputB;
input reset;
wire CTS_n_tid1_36;
wire \outB_reg[31] ;
wire \outB_reg[30] ;
wire \outB_reg[29] ;
wire \outB_reg[28] ;
wire \outB_reg[27] ;
wire \outB_reg[26] ;
wire \outB_reg[25] ;
wire \outB_reg[24] ;
wire \outB_reg[23] ;
wire \outB_reg[22] ;
wire \outB_reg[21] ;
wire \outB_reg[20] ;
wire \outB_reg[19] ;
wire \outB_reg[18] ;
wire \outB_reg[17] ;
wire \outB_reg[16] ;
wire \outB_reg[15] ;
wire \outB_reg[14] ;
wire \outB_reg[13] ;
wire \outB_reg[12] ;
wire \outB_reg[11] ;
wire \outB_reg[10] ;
wire \outB_reg[9] ;
wire \outB_reg[8] ;
wire \outB_reg[7] ;
wire \outB_reg[6] ;
wire \outB_reg[5] ;
wire \outB_reg[4] ;
wire \outB_reg[3] ;
wire \outB_reg[2] ;
wire \outB_reg[1] ;
wire \outB_reg[0] ;
wire \outA_reg[31] ;
wire \outA_reg[30] ;
wire \outA_reg[29] ;
wire \outA_reg[28] ;
wire \outA_reg[27] ;
wire \outA_reg[26] ;
wire \outA_reg[25] ;
wire \outA_reg[24] ;
wire \outA_reg[23] ;
wire \outA_reg[22] ;
wire \outA_reg[21] ;
wire \outA_reg[20] ;
wire \outA_reg[19] ;
wire \outA_reg[18] ;
wire \outA_reg[17] ;
wire \outA_reg[16] ;
wire \outA_reg[15] ;
wire \outA_reg[14] ;
wire \outA_reg[13] ;
wire \outA_reg[12] ;
wire \outA_reg[11] ;
wire \outA_reg[10] ;
wire \outA_reg[9] ;
wire \outA_reg[8] ;
wire \outA_reg[7] ;
wire \outA_reg[6] ;
wire \outA_reg[5] ;
wire \outA_reg[4] ;
wire \outA_reg[3] ;
wire \outA_reg[2] ;
wire \outA_reg[1] ;
wire \outA_reg[0] ;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire CTS_n_tid1_5;
wire CTS_n_tid1_84;
wire n_tid1_169;


registerNbits outA (.out ({result[31], result[30], result[29], result[28], result[27], 
    result[26], result[25], result[24], result[23], result[22], result[21], result[20], 
    result[19], result[18], result[17], result[16], result[15], result[14], result[13], 
    result[12], result[11], result[10], result[9], result[8], result[7], result[6], 
    result[5], result[4], result[3], result[2], result[1], result[0]}), .clk_CTS_1_PP_18 (CTS_n_tid1_84)
    , .en (en), .inp ({\outB_reg[31] , \outB_reg[30] , \outB_reg[29] , \outB_reg[28] , 
    \outB_reg[27] , \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , \outB_reg[23] , 
    \outB_reg[22] , \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , \outB_reg[18] , 
    \outB_reg[17] , \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , \outB_reg[13] , 
    \outB_reg[12] , \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , \outB_reg[8] , 
    \outB_reg[7] , \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , 
    \outB_reg[1] , \outB_reg[0] }), .reset (reset), .clk_CTS_1_PP_19 (n_tid1_169));
registerNbits__6_8 outB (.out ({result[63], result[62], result[61], result[60], result[59], 
    result[58], result[57], result[56], result[55], result[54], result[53], result[52], 
    result[51], result[50], result[49], result[48], result[47], result[46], result[45], 
    result[44], result[43], result[42], result[41], result[40], result[39], result[38], 
    result[37], result[36], result[35], result[34], result[33], result[32]}), .clk_CTS_1_PP_1 (CTS_n_tid1_5)
    , .clk_CTS_1_PP_10 (CTS_n_tid1_36), .en (en), .inp ({\outA_reg[31] , \outA_reg[30] , 
    \outA_reg[29] , \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , 
    \outA_reg[24] , \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , 
    \outA_reg[19] , \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , 
    \outA_reg[14] , \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , 
    \outA_reg[9] , \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , 
    \outA_reg[3] , \outA_reg[2] , \outA_reg[1] , \outA_reg[0] }), .reset (reset), .clk_CTS_1_PP_25 (CTS_n_tid1_84));
registerNbits__6_5 regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , 
    \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , 
    \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , 
    \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , 
    \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .en (en), .inp ({inputB[31], inputB[30], 
    inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], inputB[24], inputB[23], 
    inputB[22], inputB[21], inputB[20], inputB[19], inputB[18], inputB[17], inputB[16], 
    inputB[15], inputB[14], inputB[13], inputB[12], inputB[11], inputB[10], inputB[9], 
    inputB[8], inputB[7], inputB[6], inputB[5], inputB[4], inputB[3], inputB[2], 
    inputB[1], inputB[0]}), .reset (reset), .clk_CTS_1_PP_1 (CTS_n_tid1_5));
registerNbits__6_2 regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .en (en), .inp ({inputA[31], inputA[30], 
    inputA[29], inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], 
    inputA[22], inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], 
    inputA[15], inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], 
    inputA[8], inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], 
    inputA[1], inputA[0]}), .reset (reset), .clk_CTS_1_PP_10 (CTS_n_tid1_36));
mulTree multiplier (.out ({\outA_reg[31] , \outA_reg[30] , \outA_reg[29] , \outA_reg[28] , 
    \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , \outA_reg[24] , \outA_reg[23] , 
    \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , \outA_reg[19] , \outA_reg[18] , 
    \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , \outA_reg[14] , \outA_reg[13] , 
    \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , \outA_reg[9] , \outA_reg[8] , 
    \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , 
    \outA_reg[1] , \outA_reg[0] , \outB_reg[31] , \outB_reg[30] , \outB_reg[29] , 
    \outB_reg[28] , \outB_reg[27] , \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , 
    \outB_reg[23] , \outB_reg[22] , \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , 
    \outB_reg[18] , \outB_reg[17] , \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , 
    \outB_reg[13] , \outB_reg[12] , \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , 
    \outB_reg[8] , \outB_reg[7] , \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , 
    \outB_reg[2] , \outB_reg[1] , \outB_reg[0] }), .x ({\A_reg[31] , \A_reg[30] , 
    \A_reg[29] , \A_reg[28] , \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , 
    \A_reg[23] , \A_reg[22] , \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , 
    \A_reg[17] , \A_reg[16] , \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , 
    \A_reg[11] , \A_reg[10] , \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , 
    \A_reg[4] , \A_reg[3] , \A_reg[2] , \A_reg[1] , \A_reg[0] }), .y ({\B_reg[31] , 
    \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , \B_reg[26] , \B_reg[25] , 
    \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , \B_reg[20] , \B_reg[19] , 
    \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , \B_reg[14] , \B_reg[13] , 
    \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , 
    \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] }));
BUF_X8 CTS_L1_tid1__c1_tid1__c60 (.Z (n_tid1_169), .A (clk));

endmodule //integrationMult


