
// 	Tue Jan  3 18:08:57 2023
//	vlsi
//	localhost.localdomain

module registerNbits (clk_CTS_0_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits

module registerNbits__0_90 (clk_CTS_0_PP_8, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_8;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_25;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid0_33;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_25), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_25), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_25), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_25), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_25), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_25), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_25), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_25), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_25), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_25), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_25), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_25), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_25), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_25), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_25), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_25), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_25), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_25), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_25), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_25), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_25), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_25), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_25), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_25), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_25), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_25), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_25), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_25), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_25), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_25), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_25), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid1_25), .D (n_33));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n_tid1_25), .CK (CTS_n_tid0_33), .E (n_1), .SE (1'b0 ));
INV_X16 CTS_L6_c_tid0_24 (.ZN (CTS_n_tid0_33), .A (clk_CTS_0_PP_8));

endmodule //registerNbits__0_90

module datapath__0_74 (p_0, aux, p_1);

output [63:0] p_1;
input [63:0] aux;
input [63:0] p_0;
wire n_0;
wire n_366;
wire n_1;
wire n_365;
wire n_364;
wire n_2;
wire n_369;
wire n_363;
wire n_3;
wire n_370;
wire n_376;
wire n_372;
wire n_361;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_358;
wire n_349;
wire n_11;
wire n_5;
wire n_359;
wire n_353;
wire n_8;
wire n_356;
wire n_354;
wire n_360;
wire n_351;
wire n_347;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_344;
wire n_335;
wire n_19;
wire n_13;
wire n_345;
wire n_339;
wire n_16;
wire n_342;
wire n_340;
wire n_346;
wire n_337;
wire n_333;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_330;
wire n_321;
wire n_27;
wire n_21;
wire n_331;
wire n_325;
wire n_24;
wire n_328;
wire n_326;
wire n_332;
wire n_323;
wire n_319;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_285;
wire n_275;
wire n_35;
wire n_29;
wire n_284;
wire n_287;
wire n_277;
wire n_32;
wire n_286;
wire n_282;
wire n_279;
wire n_289;
wire n_63;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_313;
wire n_257;
wire n_43;
wire n_37;
wire n_312;
wire n_315;
wire n_259;
wire n_40;
wire n_314;
wire n_318;
wire n_261;
wire n_317;
wire n_61;
wire n_50;
wire n_49;
wire n_46;
wire n_47;
wire n_44;
wire n_296;
wire n_269;
wire n_51;
wire n_45;
wire n_295;
wire n_298;
wire n_271;
wire n_48;
wire n_297;
wire n_293;
wire n_273;
wire n_300;
wire n_59;
wire n_58;
wire n_57;
wire n_54;
wire n_55;
wire n_52;
wire n_305;
wire n_263;
wire n_65;
wire n_53;
wire n_304;
wire n_307;
wire n_266;
wire n_56;
wire n_306;
wire n_302;
wire n_267;
wire n_60;
wire n_268;
wire n_292;
wire n_62;
wire n_256;
wire n_310;
wire n_64;
wire n_274;
wire n_281;
wire n_308;
wire n_377;
wire n_373;
wire n_254;
wire n_72;
wire n_71;
wire n_68;
wire n_69;
wire n_66;
wire n_223;
wire n_213;
wire n_73;
wire n_67;
wire n_222;
wire n_225;
wire n_215;
wire n_70;
wire n_224;
wire n_220;
wire n_217;
wire n_227;
wire n_101;
wire n_80;
wire n_79;
wire n_76;
wire n_77;
wire n_74;
wire n_248;
wire n_206;
wire n_81;
wire n_75;
wire n_247;
wire n_250;
wire n_208;
wire n_78;
wire n_249;
wire n_253;
wire n_210;
wire n_252;
wire n_99;
wire n_88;
wire n_87;
wire n_84;
wire n_85;
wire n_82;
wire n_234;
wire n_192;
wire n_89;
wire n_83;
wire n_233;
wire n_236;
wire n_194;
wire n_86;
wire n_235;
wire n_231;
wire n_196;
wire n_238;
wire n_98;
wire n_97;
wire n_95;
wire n_94;
wire n_91;
wire n_90;
wire n_202;
wire n_242;
wire n_199;
wire n_103;
wire n_92;
wire n_93;
wire n_241;
wire n_200;
wire n_96;
wire n_243;
wire n_203;
wire n_204;
wire n_191;
wire n_230;
wire n_100;
wire n_205;
wire n_245;
wire n_102;
wire n_212;
wire n_219;
wire n_244;
wire n_189;
wire n_110;
wire n_109;
wire n_106;
wire n_107;
wire n_104;
wire n_186;
wire n_177;
wire n_111;
wire n_105;
wire n_187;
wire n_181;
wire n_108;
wire n_184;
wire n_182;
wire n_188;
wire n_179;
wire n_175;
wire n_118;
wire n_117;
wire n_114;
wire n_115;
wire n_112;
wire n_164;
wire n_154;
wire n_119;
wire n_113;
wire n_163;
wire n_166;
wire n_156;
wire n_116;
wire n_165;
wire n_161;
wire n_158;
wire n_168;
wire n_128;
wire n_127;
wire n_125;
wire n_124;
wire n_121;
wire n_120;
wire n_149;
wire n_172;
wire n_145;
wire n_129;
wire n_122;
wire n_123;
wire n_171;
wire n_146;
wire n_126;
wire n_173;
wire n_150;
wire n_151;
wire n_153;
wire n_160;
wire n_174;
wire n_143;
wire n_142;
wire n_140;
wire n_136;
wire n_141;
wire n_135;
wire n_131;
wire n_130;
wire n_137;
wire n_139;
wire n_133;
wire n_132;
wire n_134;
wire n_138;
wire n_379;
wire n_375;
wire n_371;
wire n_147;
wire n_144;
wire n_152;
wire n_159;
wire n_378;
wire n_374;
wire n_148;
wire n_170;
wire n_169;
wire n_155;
wire n_167;
wire n_162;
wire n_157;
wire n_176;
wire n_180;
wire n_183;
wire n_178;
wire n_185;
wire n_211;
wire n_190;
wire n_218;
wire n_197;
wire n_239;
wire n_229;
wire n_193;
wire n_237;
wire n_232;
wire n_195;
wire n_198;
wire n_201;
wire n_240;
wire n_207;
wire n_251;
wire n_246;
wire n_209;
wire n_228;
wire n_214;
wire n_226;
wire n_221;
wire n_216;
wire n_262;
wire n_255;
wire n_280;
wire n_290;
wire n_291;
wire n_301;
wire n_258;
wire n_316;
wire n_311;
wire n_260;
wire n_303;
wire n_265;
wire n_309;
wire n_264;
wire n_270;
wire n_299;
wire n_294;
wire n_272;
wire n_276;
wire n_288;
wire n_283;
wire n_278;
wire n_320;
wire n_324;
wire n_327;
wire n_322;
wire n_329;
wire n_334;
wire n_338;
wire n_341;
wire n_336;
wire n_343;
wire n_348;
wire n_352;
wire n_355;
wire n_350;
wire n_357;
wire n_362;
wire n_368;
wire n_367;


INV_X1 i_443 (.ZN (n_379), .A (p_0[61]));
INV_X1 i_442 (.ZN (n_378), .A (p_0[59]));
INV_X1 i_441 (.ZN (n_377), .A (p_0[31]));
INV_X1 i_440 (.ZN (n_376), .A (p_0[3]));
INV_X1 i_439 (.ZN (n_375), .A (aux[61]));
INV_X1 i_438 (.ZN (n_374), .A (aux[59]));
INV_X1 i_437 (.ZN (n_373), .A (aux[31]));
INV_X1 i_436 (.ZN (n_372), .A (aux[3]));
NOR2_X1 i_435 (.ZN (n_371), .A1 (p_0[60]), .A2 (aux[60]));
NAND2_X1 i_434 (.ZN (n_370), .A1 (n_376), .A2 (n_372));
NAND2_X1 i_433 (.ZN (n_369), .A1 (p_0[2]), .A2 (aux[2]));
INV_X1 i_432 (.ZN (n_368), .A (n_369));
NOR2_X1 i_431 (.ZN (n_367), .A1 (p_0[1]), .A2 (aux[1]));
NAND2_X1 i_430 (.ZN (n_366), .A1 (p_0[0]), .A2 (aux[0]));
NAND2_X1 i_429 (.ZN (n_365), .A1 (p_0[1]), .A2 (aux[1]));
AOI21_X1 i_428 (.ZN (n_364), .A (n_367), .B1 (n_366), .B2 (n_365));
OAI22_X1 i_427 (.ZN (n_363), .A1 (p_0[2]), .A2 (aux[2]), .B1 (n_368), .B2 (n_364));
OAI21_X1 i_426 (.ZN (n_362), .A (n_363), .B1 (n_376), .B2 (n_372));
NAND2_X1 i_425 (.ZN (n_361), .A1 (n_370), .A2 (n_362));
NOR2_X1 i_424 (.ZN (n_360), .A1 (p_0[7]), .A2 (aux[7]));
NOR2_X1 i_423 (.ZN (n_359), .A1 (p_0[5]), .A2 (aux[5]));
NOR2_X1 i_422 (.ZN (n_358), .A1 (p_0[6]), .A2 (aux[6]));
OR3_X1 i_421 (.ZN (n_357), .A1 (n_360), .A2 (n_358), .A3 (n_359));
NOR2_X1 i_420 (.ZN (n_356), .A1 (p_0[4]), .A2 (aux[4]));
NOR3_X1 i_419 (.ZN (n_355), .A1 (n_357), .A2 (n_356), .A3 (n_361));
NAND2_X1 i_418 (.ZN (n_354), .A1 (p_0[4]), .A2 (aux[4]));
NAND2_X1 i_417 (.ZN (n_353), .A1 (p_0[5]), .A2 (aux[5]));
AOI21_X1 i_416 (.ZN (n_352), .A (n_357), .B1 (n_354), .B2 (n_353));
AND2_X1 i_415 (.ZN (n_351), .A1 (p_0[7]), .A2 (aux[7]));
NAND2_X1 i_414 (.ZN (n_350), .A1 (p_0[6]), .A2 (aux[6]));
INV_X1 i_413 (.ZN (n_349), .A (n_350));
NOR2_X1 i_412 (.ZN (n_348), .A1 (n_360), .A2 (n_350));
NOR4_X1 i_411 (.ZN (n_347), .A1 (n_351), .A2 (n_348), .A3 (n_352), .A4 (n_355));
NOR2_X1 i_410 (.ZN (n_346), .A1 (p_0[11]), .A2 (aux[11]));
NOR2_X1 i_409 (.ZN (n_345), .A1 (p_0[9]), .A2 (aux[9]));
NOR2_X1 i_408 (.ZN (n_344), .A1 (p_0[10]), .A2 (aux[10]));
OR3_X1 i_407 (.ZN (n_343), .A1 (n_346), .A2 (n_344), .A3 (n_345));
NOR2_X1 i_406 (.ZN (n_342), .A1 (p_0[8]), .A2 (aux[8]));
NOR3_X1 i_405 (.ZN (n_341), .A1 (n_343), .A2 (n_342), .A3 (n_347));
NAND2_X1 i_404 (.ZN (n_340), .A1 (p_0[8]), .A2 (aux[8]));
NAND2_X1 i_403 (.ZN (n_339), .A1 (p_0[9]), .A2 (aux[9]));
AOI21_X1 i_402 (.ZN (n_338), .A (n_343), .B1 (n_340), .B2 (n_339));
AND2_X1 i_401 (.ZN (n_337), .A1 (p_0[11]), .A2 (aux[11]));
NAND2_X1 i_400 (.ZN (n_336), .A1 (p_0[10]), .A2 (aux[10]));
INV_X1 i_399 (.ZN (n_335), .A (n_336));
NOR2_X1 i_398 (.ZN (n_334), .A1 (n_346), .A2 (n_336));
NOR4_X1 i_397 (.ZN (n_333), .A1 (n_337), .A2 (n_334), .A3 (n_338), .A4 (n_341));
NOR2_X1 i_396 (.ZN (n_332), .A1 (p_0[15]), .A2 (aux[15]));
NOR2_X1 i_395 (.ZN (n_331), .A1 (p_0[13]), .A2 (aux[13]));
NOR2_X1 i_394 (.ZN (n_330), .A1 (p_0[14]), .A2 (aux[14]));
OR3_X1 i_393 (.ZN (n_329), .A1 (n_332), .A2 (n_330), .A3 (n_331));
NOR2_X1 i_392 (.ZN (n_328), .A1 (p_0[12]), .A2 (aux[12]));
NOR3_X1 i_391 (.ZN (n_327), .A1 (n_329), .A2 (n_328), .A3 (n_333));
NAND2_X1 i_390 (.ZN (n_326), .A1 (p_0[12]), .A2 (aux[12]));
NAND2_X1 i_389 (.ZN (n_325), .A1 (p_0[13]), .A2 (aux[13]));
AOI21_X1 i_388 (.ZN (n_324), .A (n_329), .B1 (n_326), .B2 (n_325));
AND2_X1 i_387 (.ZN (n_323), .A1 (p_0[15]), .A2 (aux[15]));
NAND2_X1 i_386 (.ZN (n_322), .A1 (p_0[14]), .A2 (aux[14]));
INV_X1 i_385 (.ZN (n_321), .A (n_322));
NOR2_X1 i_384 (.ZN (n_320), .A1 (n_332), .A2 (n_322));
NOR4_X2 i_383 (.ZN (n_319), .A1 (n_323), .A2 (n_320), .A3 (n_324), .A4 (n_327));
NOR2_X1 i_382 (.ZN (n_318), .A1 (p_0[20]), .A2 (aux[20]));
NOR2_X1 i_381 (.ZN (n_317), .A1 (p_0[23]), .A2 (aux[23]));
INV_X1 i_380 (.ZN (n_316), .A (n_317));
NOR2_X1 i_379 (.ZN (n_315), .A1 (p_0[21]), .A2 (aux[21]));
INV_X1 i_378 (.ZN (n_314), .A (n_315));
NOR2_X1 i_377 (.ZN (n_313), .A1 (p_0[22]), .A2 (aux[22]));
INV_X1 i_376 (.ZN (n_312), .A (n_313));
NAND3_X1 i_375 (.ZN (n_311), .A1 (n_316), .A2 (n_312), .A3 (n_314));
OR2_X1 i_374 (.ZN (n_310), .A1 (n_318), .A2 (n_311));
NOR2_X1 i_373 (.ZN (n_309), .A1 (p_0[31]), .A2 (aux[31]));
INV_X1 i_372 (.ZN (n_308), .A (n_309));
NOR2_X1 i_371 (.ZN (n_307), .A1 (p_0[29]), .A2 (aux[29]));
INV_X1 i_370 (.ZN (n_306), .A (n_307));
NOR2_X1 i_369 (.ZN (n_305), .A1 (p_0[30]), .A2 (aux[30]));
INV_X1 i_368 (.ZN (n_304), .A (n_305));
NAND3_X1 i_367 (.ZN (n_303), .A1 (n_308), .A2 (n_304), .A3 (n_306));
NOR2_X1 i_366 (.ZN (n_302), .A1 (p_0[28]), .A2 (aux[28]));
OR2_X1 i_365 (.ZN (n_301), .A1 (n_303), .A2 (n_302));
NOR2_X1 i_364 (.ZN (n_300), .A1 (p_0[27]), .A2 (aux[27]));
INV_X1 i_363 (.ZN (n_299), .A (n_300));
NOR2_X1 i_362 (.ZN (n_298), .A1 (p_0[25]), .A2 (aux[25]));
INV_X1 i_361 (.ZN (n_297), .A (n_298));
NOR2_X1 i_360 (.ZN (n_296), .A1 (p_0[26]), .A2 (aux[26]));
INV_X1 i_359 (.ZN (n_295), .A (n_296));
NAND3_X1 i_358 (.ZN (n_294), .A1 (n_299), .A2 (n_295), .A3 (n_297));
NOR2_X1 i_357 (.ZN (n_293), .A1 (p_0[24]), .A2 (aux[24]));
OR2_X1 i_356 (.ZN (n_292), .A1 (n_294), .A2 (n_293));
OR2_X1 i_355 (.ZN (n_291), .A1 (n_301), .A2 (n_292));
OR2_X1 i_354 (.ZN (n_290), .A1 (n_310), .A2 (n_291));
NOR2_X1 i_353 (.ZN (n_289), .A1 (p_0[19]), .A2 (aux[19]));
INV_X1 i_352 (.ZN (n_288), .A (n_289));
NOR2_X1 i_351 (.ZN (n_287), .A1 (p_0[17]), .A2 (aux[17]));
INV_X1 i_350 (.ZN (n_286), .A (n_287));
NOR2_X1 i_349 (.ZN (n_285), .A1 (p_0[18]), .A2 (aux[18]));
INV_X1 i_348 (.ZN (n_284), .A (n_285));
NAND3_X1 i_347 (.ZN (n_283), .A1 (n_288), .A2 (n_284), .A3 (n_286));
NOR2_X1 i_346 (.ZN (n_282), .A1 (p_0[16]), .A2 (aux[16]));
OR2_X1 i_345 (.ZN (n_281), .A1 (n_283), .A2 (n_282));
NOR3_X1 i_344 (.ZN (n_280), .A1 (n_290), .A2 (n_281), .A3 (n_319));
NAND2_X1 i_343 (.ZN (n_279), .A1 (p_0[16]), .A2 (aux[16]));
NAND2_X1 i_342 (.ZN (n_278), .A1 (p_0[17]), .A2 (aux[17]));
INV_X1 i_341 (.ZN (n_277), .A (n_278));
AOI21_X1 i_340 (.ZN (n_276), .A (n_283), .B1 (n_279), .B2 (n_278));
AND2_X1 i_339 (.ZN (n_275), .A1 (p_0[18]), .A2 (aux[18]));
AOI221_X1 i_338 (.ZN (n_274), .A (n_276), .B1 (p_0[19]), .B2 (aux[19]), .C1 (n_288), .C2 (n_275));
NAND2_X1 i_337 (.ZN (n_273), .A1 (p_0[24]), .A2 (aux[24]));
NAND2_X1 i_336 (.ZN (n_272), .A1 (p_0[25]), .A2 (aux[25]));
INV_X1 i_335 (.ZN (n_271), .A (n_272));
AOI21_X1 i_334 (.ZN (n_270), .A (n_294), .B1 (n_273), .B2 (n_272));
AND2_X1 i_333 (.ZN (n_269), .A1 (p_0[26]), .A2 (aux[26]));
AOI221_X1 i_332 (.ZN (n_268), .A (n_270), .B1 (p_0[27]), .B2 (aux[27]), .C1 (n_299), .C2 (n_269));
NAND2_X1 i_331 (.ZN (n_267), .A1 (p_0[28]), .A2 (aux[28]));
AND2_X1 i_330 (.ZN (n_266), .A1 (p_0[29]), .A2 (aux[29]));
AOI21_X1 i_329 (.ZN (n_265), .A (n_266), .B1 (p_0[28]), .B2 (aux[28]));
NAND2_X1 i_328 (.ZN (n_264), .A1 (p_0[30]), .A2 (aux[30]));
INV_X1 i_327 (.ZN (n_263), .A (n_264));
OAI222_X1 i_326 (.ZN (n_262), .A1 (n_303), .A2 (n_265), .B1 (n_309), .B2 (n_264), .C1 (n_377), .C2 (n_373));
NAND2_X1 i_325 (.ZN (n_261), .A1 (p_0[20]), .A2 (aux[20]));
NAND2_X1 i_324 (.ZN (n_260), .A1 (p_0[21]), .A2 (aux[21]));
INV_X1 i_323 (.ZN (n_259), .A (n_260));
AOI21_X1 i_322 (.ZN (n_258), .A (n_311), .B1 (n_261), .B2 (n_260));
AND2_X1 i_321 (.ZN (n_257), .A1 (p_0[22]), .A2 (aux[22]));
AOI221_X1 i_320 (.ZN (n_256), .A (n_258), .B1 (p_0[23]), .B2 (aux[23]), .C1 (n_316), .C2 (n_257));
OAI222_X1 i_319 (.ZN (n_255), .A1 (n_290), .A2 (n_274), .B1 (n_291), .B2 (n_256), .C1 (n_301), .C2 (n_268));
NOR3_X2 i_318 (.ZN (n_254), .A1 (n_262), .A2 (n_255), .A3 (n_280));
NOR2_X1 i_317 (.ZN (n_253), .A1 (p_0[36]), .A2 (aux[36]));
NOR2_X1 i_316 (.ZN (n_252), .A1 (p_0[39]), .A2 (aux[39]));
INV_X1 i_315 (.ZN (n_251), .A (n_252));
NOR2_X1 i_314 (.ZN (n_250), .A1 (p_0[37]), .A2 (aux[37]));
INV_X1 i_313 (.ZN (n_249), .A (n_250));
NOR2_X1 i_312 (.ZN (n_248), .A1 (p_0[38]), .A2 (aux[38]));
INV_X1 i_311 (.ZN (n_247), .A (n_248));
NAND3_X1 i_310 (.ZN (n_246), .A1 (n_251), .A2 (n_247), .A3 (n_249));
OR2_X1 i_309 (.ZN (n_245), .A1 (n_253), .A2 (n_246));
NOR2_X1 i_308 (.ZN (n_244), .A1 (p_0[47]), .A2 (aux[47]));
NOR2_X1 i_307 (.ZN (n_243), .A1 (p_0[45]), .A2 (aux[45]));
NOR2_X1 i_306 (.ZN (n_242), .A1 (p_0[46]), .A2 (aux[46]));
NOR2_X1 i_305 (.ZN (n_241), .A1 (n_243), .A2 (n_242));
NOR3_X1 i_304 (.ZN (n_240), .A1 (n_244), .A2 (n_242), .A3 (n_243));
OAI21_X1 i_303 (.ZN (n_239), .A (n_240), .B1 (p_0[44]), .B2 (aux[44]));
NOR2_X1 i_302 (.ZN (n_238), .A1 (p_0[43]), .A2 (aux[43]));
INV_X1 i_301 (.ZN (n_237), .A (n_238));
NOR2_X1 i_300 (.ZN (n_236), .A1 (p_0[41]), .A2 (aux[41]));
INV_X1 i_299 (.ZN (n_235), .A (n_236));
NOR2_X1 i_298 (.ZN (n_234), .A1 (p_0[42]), .A2 (aux[42]));
INV_X1 i_297 (.ZN (n_233), .A (n_234));
NAND3_X1 i_296 (.ZN (n_232), .A1 (n_237), .A2 (n_233), .A3 (n_235));
NOR2_X1 i_295 (.ZN (n_231), .A1 (p_0[40]), .A2 (aux[40]));
OR2_X1 i_294 (.ZN (n_230), .A1 (n_232), .A2 (n_231));
OR2_X1 i_293 (.ZN (n_229), .A1 (n_239), .A2 (n_230));
OR2_X1 i_292 (.ZN (n_228), .A1 (n_245), .A2 (n_229));
NOR2_X1 i_291 (.ZN (n_227), .A1 (p_0[35]), .A2 (aux[35]));
INV_X1 i_290 (.ZN (n_226), .A (n_227));
NOR2_X1 i_289 (.ZN (n_225), .A1 (p_0[33]), .A2 (aux[33]));
INV_X1 i_288 (.ZN (n_224), .A (n_225));
NOR2_X1 i_287 (.ZN (n_223), .A1 (p_0[34]), .A2 (aux[34]));
INV_X1 i_286 (.ZN (n_222), .A (n_223));
NAND3_X1 i_285 (.ZN (n_221), .A1 (n_226), .A2 (n_222), .A3 (n_224));
NOR2_X1 i_284 (.ZN (n_220), .A1 (p_0[32]), .A2 (aux[32]));
OR2_X1 i_283 (.ZN (n_219), .A1 (n_221), .A2 (n_220));
NOR3_X1 i_282 (.ZN (n_218), .A1 (n_228), .A2 (n_219), .A3 (n_254));
NAND2_X1 i_281 (.ZN (n_217), .A1 (p_0[32]), .A2 (aux[32]));
NAND2_X1 i_280 (.ZN (n_216), .A1 (p_0[33]), .A2 (aux[33]));
INV_X1 i_279 (.ZN (n_215), .A (n_216));
AOI21_X1 i_278 (.ZN (n_214), .A (n_221), .B1 (n_217), .B2 (n_216));
AND2_X1 i_277 (.ZN (n_213), .A1 (p_0[34]), .A2 (aux[34]));
AOI221_X1 i_276 (.ZN (n_212), .A (n_214), .B1 (p_0[35]), .B2 (aux[35]), .C1 (n_226), .C2 (n_213));
NOR2_X1 i_275 (.ZN (n_211), .A1 (n_228), .A2 (n_212));
NAND2_X1 i_274 (.ZN (n_210), .A1 (p_0[36]), .A2 (aux[36]));
NAND2_X1 i_273 (.ZN (n_209), .A1 (p_0[37]), .A2 (aux[37]));
INV_X1 i_272 (.ZN (n_208), .A (n_209));
AOI21_X1 i_271 (.ZN (n_207), .A (n_246), .B1 (n_210), .B2 (n_209));
AND2_X1 i_270 (.ZN (n_206), .A1 (p_0[38]), .A2 (aux[38]));
AOI221_X1 i_269 (.ZN (n_205), .A (n_207), .B1 (p_0[39]), .B2 (aux[39]), .C1 (n_251), .C2 (n_206));
NAND2_X1 i_268 (.ZN (n_204), .A1 (p_0[44]), .A2 (aux[44]));
INV_X1 i_267 (.ZN (n_203), .A (n_204));
AND2_X1 i_266 (.ZN (n_202), .A1 (p_0[45]), .A2 (aux[45]));
OAI21_X1 i_265 (.ZN (n_201), .A (n_240), .B1 (n_203), .B2 (n_202));
NAND2_X1 i_264 (.ZN (n_200), .A1 (p_0[46]), .A2 (aux[46]));
INV_X1 i_263 (.ZN (n_199), .A (n_200));
OAI21_X1 i_262 (.ZN (n_198), .A (n_201), .B1 (n_244), .B2 (n_200));
AOI21_X1 i_261 (.ZN (n_197), .A (n_198), .B1 (p_0[47]), .B2 (aux[47]));
NAND2_X1 i_260 (.ZN (n_196), .A1 (p_0[40]), .A2 (aux[40]));
NAND2_X1 i_259 (.ZN (n_195), .A1 (p_0[41]), .A2 (aux[41]));
INV_X1 i_258 (.ZN (n_194), .A (n_195));
AOI21_X1 i_257 (.ZN (n_193), .A (n_232), .B1 (n_196), .B2 (n_195));
AND2_X1 i_256 (.ZN (n_192), .A1 (p_0[42]), .A2 (aux[42]));
AOI221_X1 i_255 (.ZN (n_191), .A (n_193), .B1 (p_0[43]), .B2 (aux[43]), .C1 (n_237), .C2 (n_192));
OAI221_X1 i_254 (.ZN (n_190), .A (n_197), .B1 (n_239), .B2 (n_191), .C1 (n_229), .C2 (n_205));
NOR3_X1 i_253 (.ZN (n_189), .A1 (n_211), .A2 (n_190), .A3 (n_218));
NOR2_X1 i_252 (.ZN (n_188), .A1 (p_0[51]), .A2 (aux[51]));
NOR2_X1 i_251 (.ZN (n_187), .A1 (p_0[49]), .A2 (aux[49]));
NOR2_X1 i_250 (.ZN (n_186), .A1 (p_0[50]), .A2 (aux[50]));
OR3_X1 i_249 (.ZN (n_185), .A1 (n_188), .A2 (n_186), .A3 (n_187));
NOR2_X1 i_248 (.ZN (n_184), .A1 (p_0[48]), .A2 (aux[48]));
NOR3_X1 i_247 (.ZN (n_183), .A1 (n_185), .A2 (n_184), .A3 (n_189));
NAND2_X1 i_246 (.ZN (n_182), .A1 (p_0[48]), .A2 (aux[48]));
NAND2_X1 i_245 (.ZN (n_181), .A1 (p_0[49]), .A2 (aux[49]));
AOI21_X1 i_244 (.ZN (n_180), .A (n_185), .B1 (n_182), .B2 (n_181));
AND2_X1 i_243 (.ZN (n_179), .A1 (p_0[51]), .A2 (aux[51]));
NAND2_X1 i_242 (.ZN (n_178), .A1 (p_0[50]), .A2 (aux[50]));
INV_X1 i_241 (.ZN (n_177), .A (n_178));
NOR2_X1 i_240 (.ZN (n_176), .A1 (n_188), .A2 (n_178));
NOR4_X2 i_239 (.ZN (n_175), .A1 (n_179), .A2 (n_176), .A3 (n_180), .A4 (n_183));
NOR2_X1 i_238 (.ZN (n_174), .A1 (p_0[59]), .A2 (aux[59]));
NOR2_X1 i_237 (.ZN (n_173), .A1 (p_0[57]), .A2 (aux[57]));
NOR2_X1 i_236 (.ZN (n_172), .A1 (p_0[58]), .A2 (aux[58]));
NOR2_X1 i_235 (.ZN (n_171), .A1 (n_173), .A2 (n_172));
NOR3_X1 i_234 (.ZN (n_170), .A1 (n_174), .A2 (n_172), .A3 (n_173));
OAI21_X1 i_233 (.ZN (n_169), .A (n_170), .B1 (p_0[56]), .B2 (aux[56]));
NOR2_X1 i_232 (.ZN (n_168), .A1 (p_0[55]), .A2 (aux[55]));
INV_X1 i_231 (.ZN (n_167), .A (n_168));
NOR2_X1 i_230 (.ZN (n_166), .A1 (p_0[53]), .A2 (aux[53]));
INV_X1 i_229 (.ZN (n_165), .A (n_166));
NOR2_X1 i_228 (.ZN (n_164), .A1 (p_0[54]), .A2 (aux[54]));
INV_X1 i_227 (.ZN (n_163), .A (n_164));
NAND3_X1 i_226 (.ZN (n_162), .A1 (n_167), .A2 (n_163), .A3 (n_165));
NOR2_X1 i_225 (.ZN (n_161), .A1 (p_0[52]), .A2 (aux[52]));
OR2_X1 i_224 (.ZN (n_160), .A1 (n_162), .A2 (n_161));
NOR3_X1 i_223 (.ZN (n_159), .A1 (n_169), .A2 (n_160), .A3 (n_175));
NAND2_X1 i_222 (.ZN (n_158), .A1 (p_0[52]), .A2 (aux[52]));
NAND2_X1 i_221 (.ZN (n_157), .A1 (p_0[53]), .A2 (aux[53]));
INV_X1 i_220 (.ZN (n_156), .A (n_157));
AOI21_X1 i_219 (.ZN (n_155), .A (n_162), .B1 (n_158), .B2 (n_157));
AND2_X1 i_218 (.ZN (n_154), .A1 (p_0[54]), .A2 (aux[54]));
AOI221_X1 i_217 (.ZN (n_153), .A (n_155), .B1 (p_0[55]), .B2 (aux[55]), .C1 (n_167), .C2 (n_154));
NOR2_X1 i_216 (.ZN (n_152), .A1 (n_169), .A2 (n_153));
NAND2_X1 i_215 (.ZN (n_151), .A1 (p_0[56]), .A2 (aux[56]));
INV_X1 i_214 (.ZN (n_150), .A (n_151));
AND2_X1 i_213 (.ZN (n_149), .A1 (p_0[57]), .A2 (aux[57]));
OAI21_X1 i_212 (.ZN (n_148), .A (n_170), .B1 (n_150), .B2 (n_149));
INV_X1 i_211 (.ZN (n_147), .A (n_148));
NAND2_X1 i_210 (.ZN (n_146), .A1 (p_0[58]), .A2 (aux[58]));
INV_X1 i_209 (.ZN (n_145), .A (n_146));
OAI22_X1 i_208 (.ZN (n_144), .A1 (n_378), .A2 (n_374), .B1 (n_174), .B2 (n_146));
NOR4_X1 i_207 (.ZN (n_143), .A1 (n_147), .A2 (n_144), .A3 (n_152), .A4 (n_159));
AOI21_X1 i_206 (.ZN (n_142), .A (n_371), .B1 (p_0[60]), .B2 (aux[60]));
AOI21_X1 i_205 (.ZN (n_141), .A (n_371), .B1 (n_143), .B2 (n_142));
INV_X1 i_204 (.ZN (n_140), .A (n_141));
NAND2_X1 i_203 (.ZN (n_139), .A1 (p_0[62]), .A2 (aux[62]));
INV_X1 i_202 (.ZN (n_138), .A (n_139));
NAND2_X1 i_201 (.ZN (n_137), .A1 (n_379), .A2 (n_375));
OAI21_X1 i_200 (.ZN (n_136), .A (n_137), .B1 (n_379), .B2 (n_375));
INV_X1 i_199 (.ZN (n_135), .A (n_136));
NAND3_X1 i_198 (.ZN (n_134), .A1 (n_139), .A2 (n_135), .A3 (n_140));
OAI221_X1 i_197 (.ZN (n_133), .A (n_134), .B1 (p_0[62]), .B2 (aux[62]), .C1 (n_138), .C2 (n_137));
XNOR2_X1 i_196 (.ZN (n_132), .A (p_0[63]), .B (aux[63]));
XOR2_X1 i_195 (.Z (p_1[63]), .A (n_133), .B (n_132));
OAI21_X1 i_194 (.ZN (n_131), .A (n_139), .B1 (p_0[62]), .B2 (aux[62]));
AOI22_X1 i_193 (.ZN (n_130), .A1 (p_0[61]), .A2 (aux[61]), .B1 (n_141), .B2 (n_137));
XOR2_X1 i_192 (.Z (p_1[62]), .A (n_131), .B (n_130));
AOI22_X1 i_191 (.ZN (p_1[61]), .A1 (n_140), .A2 (n_136), .B1 (n_141), .B2 (n_135));
XNOR2_X1 i_190 (.ZN (p_1[60]), .A (n_143), .B (n_142));
AOI21_X1 i_189 (.ZN (n_129), .A (n_174), .B1 (p_0[59]), .B2 (aux[59]));
OAI21_X1 i_188 (.ZN (n_128), .A (n_153), .B1 (n_175), .B2 (n_160));
OAI21_X1 i_187 (.ZN (n_127), .A (n_151), .B1 (p_0[56]), .B2 (aux[56]));
OAI22_X1 i_186 (.ZN (n_126), .A1 (p_0[56]), .A2 (aux[56]), .B1 (n_150), .B2 (n_128));
INV_X1 i_185 (.ZN (n_125), .A (n_126));
NOR2_X1 i_184 (.ZN (n_124), .A1 (n_173), .A2 (n_149));
NAND3_X1 i_183 (.ZN (n_123), .A1 (n_146), .A2 (n_124), .A3 (n_126));
OAI21_X1 i_182 (.ZN (n_122), .A (n_123), .B1 (n_171), .B2 (n_145));
XNOR2_X1 i_181 (.ZN (p_1[59]), .A (n_129), .B (n_122));
NOR2_X1 i_180 (.ZN (n_121), .A1 (n_172), .A2 (n_145));
OAI22_X1 i_179 (.ZN (n_120), .A1 (p_0[57]), .A2 (aux[57]), .B1 (n_149), .B2 (n_125));
XNOR2_X1 i_178 (.ZN (p_1[58]), .A (n_121), .B (n_120));
XOR2_X1 i_177 (.Z (p_1[57]), .A (n_125), .B (n_124));
XNOR2_X1 i_176 (.ZN (p_1[56]), .A (n_128), .B (n_127));
AOI21_X1 i_175 (.ZN (n_119), .A (n_168), .B1 (p_0[55]), .B2 (aux[55]));
OAI21_X1 i_174 (.ZN (n_118), .A (n_158), .B1 (p_0[52]), .B2 (aux[52]));
AOI21_X1 i_173 (.ZN (n_117), .A (n_161), .B1 (n_175), .B2 (n_158));
OAI21_X1 i_172 (.ZN (n_116), .A (n_165), .B1 (n_156), .B2 (n_117));
INV_X1 i_171 (.ZN (n_115), .A (n_116));
NOR2_X1 i_170 (.ZN (n_114), .A1 (n_166), .A2 (n_156));
OAI21_X1 i_169 (.ZN (n_113), .A (n_163), .B1 (n_154), .B2 (n_115));
XNOR2_X1 i_168 (.ZN (p_1[55]), .A (n_119), .B (n_113));
NOR2_X1 i_167 (.ZN (n_112), .A1 (n_164), .A2 (n_154));
XOR2_X1 i_166 (.Z (p_1[54]), .A (n_115), .B (n_112));
XOR2_X1 i_165 (.Z (p_1[53]), .A (n_117), .B (n_114));
XOR2_X1 i_164 (.Z (p_1[52]), .A (n_175), .B (n_118));
NOR2_X1 i_163 (.ZN (n_111), .A1 (n_188), .A2 (n_179));
OAI21_X1 i_162 (.ZN (n_110), .A (n_182), .B1 (p_0[48]), .B2 (aux[48]));
AOI21_X1 i_161 (.ZN (n_109), .A (n_184), .B1 (n_189), .B2 (n_182));
INV_X1 i_160 (.ZN (n_108), .A (n_109));
AOI21_X1 i_159 (.ZN (n_107), .A (n_187), .B1 (n_181), .B2 (n_108));
AOI21_X1 i_158 (.ZN (n_106), .A (n_187), .B1 (p_0[49]), .B2 (aux[49]));
OAI22_X1 i_157 (.ZN (n_105), .A1 (p_0[50]), .A2 (aux[50]), .B1 (n_177), .B2 (n_107));
XNOR2_X1 i_156 (.ZN (p_1[51]), .A (n_111), .B (n_105));
NOR2_X1 i_155 (.ZN (n_104), .A1 (n_186), .A2 (n_177));
XOR2_X1 i_154 (.Z (p_1[50]), .A (n_107), .B (n_104));
XOR2_X1 i_153 (.Z (p_1[49]), .A (n_109), .B (n_106));
XOR2_X1 i_152 (.Z (p_1[48]), .A (n_189), .B (n_110));
AOI21_X1 i_151 (.ZN (n_103), .A (n_244), .B1 (p_0[47]), .B2 (aux[47]));
OAI21_X1 i_150 (.ZN (n_102), .A (n_212), .B1 (n_254), .B2 (n_219));
INV_X1 i_149 (.ZN (n_101), .A (n_102));
OAI21_X1 i_148 (.ZN (n_100), .A (n_205), .B1 (n_245), .B2 (n_101));
INV_X1 i_147 (.ZN (n_99), .A (n_100));
OAI21_X1 i_146 (.ZN (n_98), .A (n_191), .B1 (n_230), .B2 (n_99));
OAI21_X1 i_145 (.ZN (n_97), .A (n_204), .B1 (p_0[44]), .B2 (aux[44]));
OAI22_X1 i_144 (.ZN (n_96), .A1 (p_0[44]), .A2 (aux[44]), .B1 (n_203), .B2 (n_98));
INV_X1 i_143 (.ZN (n_95), .A (n_96));
NOR2_X1 i_142 (.ZN (n_94), .A1 (n_243), .A2 (n_202));
NAND3_X1 i_141 (.ZN (n_93), .A1 (n_200), .A2 (n_94), .A3 (n_96));
OAI21_X1 i_140 (.ZN (n_92), .A (n_93), .B1 (n_241), .B2 (n_199));
XNOR2_X1 i_139 (.ZN (p_1[47]), .A (n_103), .B (n_92));
NOR2_X1 i_138 (.ZN (n_91), .A1 (n_242), .A2 (n_199));
OAI22_X1 i_137 (.ZN (n_90), .A1 (p_0[45]), .A2 (aux[45]), .B1 (n_202), .B2 (n_95));
XNOR2_X1 i_136 (.ZN (p_1[46]), .A (n_91), .B (n_90));
XOR2_X1 i_135 (.Z (p_1[45]), .A (n_95), .B (n_94));
XNOR2_X1 i_134 (.ZN (p_1[44]), .A (n_98), .B (n_97));
AOI21_X1 i_133 (.ZN (n_89), .A (n_238), .B1 (p_0[43]), .B2 (aux[43]));
OAI21_X1 i_132 (.ZN (n_88), .A (n_196), .B1 (p_0[40]), .B2 (aux[40]));
AOI21_X1 i_131 (.ZN (n_87), .A (n_231), .B1 (n_196), .B2 (n_99));
OAI21_X1 i_130 (.ZN (n_86), .A (n_235), .B1 (n_194), .B2 (n_87));
INV_X1 i_129 (.ZN (n_85), .A (n_86));
NOR2_X1 i_128 (.ZN (n_84), .A1 (n_236), .A2 (n_194));
OAI21_X1 i_127 (.ZN (n_83), .A (n_233), .B1 (n_192), .B2 (n_85));
XNOR2_X1 i_126 (.ZN (p_1[43]), .A (n_89), .B (n_83));
NOR2_X1 i_125 (.ZN (n_82), .A1 (n_234), .A2 (n_192));
XOR2_X1 i_124 (.Z (p_1[42]), .A (n_85), .B (n_82));
XOR2_X1 i_123 (.Z (p_1[41]), .A (n_87), .B (n_84));
XOR2_X1 i_122 (.Z (p_1[40]), .A (n_99), .B (n_88));
AOI21_X1 i_121 (.ZN (n_81), .A (n_252), .B1 (p_0[39]), .B2 (aux[39]));
OAI21_X1 i_120 (.ZN (n_80), .A (n_210), .B1 (p_0[36]), .B2 (aux[36]));
AOI21_X1 i_119 (.ZN (n_79), .A (n_253), .B1 (n_210), .B2 (n_101));
OAI21_X1 i_118 (.ZN (n_78), .A (n_249), .B1 (n_208), .B2 (n_79));
INV_X1 i_117 (.ZN (n_77), .A (n_78));
NOR2_X1 i_116 (.ZN (n_76), .A1 (n_250), .A2 (n_208));
OAI21_X1 i_115 (.ZN (n_75), .A (n_247), .B1 (n_206), .B2 (n_77));
XNOR2_X1 i_114 (.ZN (p_1[39]), .A (n_81), .B (n_75));
NOR2_X1 i_113 (.ZN (n_74), .A1 (n_248), .A2 (n_206));
XOR2_X1 i_112 (.Z (p_1[38]), .A (n_77), .B (n_74));
XOR2_X1 i_111 (.Z (p_1[37]), .A (n_79), .B (n_76));
XOR2_X1 i_110 (.Z (p_1[36]), .A (n_101), .B (n_80));
AOI21_X1 i_109 (.ZN (n_73), .A (n_227), .B1 (p_0[35]), .B2 (aux[35]));
OAI21_X1 i_108 (.ZN (n_72), .A (n_217), .B1 (p_0[32]), .B2 (aux[32]));
AOI21_X1 i_107 (.ZN (n_71), .A (n_220), .B1 (n_254), .B2 (n_217));
OAI21_X1 i_106 (.ZN (n_70), .A (n_224), .B1 (n_215), .B2 (n_71));
INV_X1 i_105 (.ZN (n_69), .A (n_70));
NOR2_X1 i_104 (.ZN (n_68), .A1 (n_225), .A2 (n_215));
OAI21_X1 i_103 (.ZN (n_67), .A (n_222), .B1 (n_213), .B2 (n_69));
XNOR2_X1 i_102 (.ZN (p_1[35]), .A (n_73), .B (n_67));
NOR2_X1 i_101 (.ZN (n_66), .A1 (n_223), .A2 (n_213));
XOR2_X1 i_100 (.Z (p_1[34]), .A (n_69), .B (n_66));
XOR2_X1 i_99 (.Z (p_1[33]), .A (n_71), .B (n_68));
XOR2_X1 i_98 (.Z (p_1[32]), .A (n_254), .B (n_72));
OAI21_X1 i_97 (.ZN (n_65), .A (n_308), .B1 (n_377), .B2 (n_373));
OAI21_X1 i_96 (.ZN (n_64), .A (n_274), .B1 (n_319), .B2 (n_281));
INV_X1 i_95 (.ZN (n_63), .A (n_64));
OAI21_X1 i_94 (.ZN (n_62), .A (n_256), .B1 (n_310), .B2 (n_63));
INV_X1 i_93 (.ZN (n_61), .A (n_62));
OAI21_X1 i_92 (.ZN (n_60), .A (n_268), .B1 (n_292), .B2 (n_61));
INV_X1 i_91 (.ZN (n_59), .A (n_60));
OAI21_X1 i_90 (.ZN (n_58), .A (n_267), .B1 (p_0[28]), .B2 (aux[28]));
AOI21_X1 i_89 (.ZN (n_57), .A (n_302), .B1 (n_267), .B2 (n_59));
OAI21_X1 i_88 (.ZN (n_56), .A (n_306), .B1 (n_266), .B2 (n_57));
INV_X1 i_87 (.ZN (n_55), .A (n_56));
NOR2_X1 i_86 (.ZN (n_54), .A1 (n_307), .A2 (n_266));
OAI21_X1 i_85 (.ZN (n_53), .A (n_304), .B1 (n_263), .B2 (n_55));
XOR2_X1 i_84 (.Z (p_1[31]), .A (n_65), .B (n_53));
NOR2_X1 i_83 (.ZN (n_52), .A1 (n_305), .A2 (n_263));
XOR2_X1 i_82 (.Z (p_1[30]), .A (n_55), .B (n_52));
XOR2_X1 i_81 (.Z (p_1[29]), .A (n_57), .B (n_54));
XOR2_X1 i_80 (.Z (p_1[28]), .A (n_59), .B (n_58));
AOI21_X1 i_79 (.ZN (n_51), .A (n_300), .B1 (p_0[27]), .B2 (aux[27]));
OAI21_X1 i_78 (.ZN (n_50), .A (n_273), .B1 (p_0[24]), .B2 (aux[24]));
AOI21_X1 i_77 (.ZN (n_49), .A (n_293), .B1 (n_273), .B2 (n_61));
OAI21_X1 i_76 (.ZN (n_48), .A (n_297), .B1 (n_271), .B2 (n_49));
INV_X1 i_75 (.ZN (n_47), .A (n_48));
NOR2_X1 i_74 (.ZN (n_46), .A1 (n_298), .A2 (n_271));
OAI21_X1 i_73 (.ZN (n_45), .A (n_295), .B1 (n_269), .B2 (n_47));
XNOR2_X1 i_72 (.ZN (p_1[27]), .A (n_51), .B (n_45));
NOR2_X1 i_71 (.ZN (n_44), .A1 (n_296), .A2 (n_269));
XOR2_X1 i_70 (.Z (p_1[26]), .A (n_47), .B (n_44));
XOR2_X1 i_69 (.Z (p_1[25]), .A (n_49), .B (n_46));
XOR2_X1 i_68 (.Z (p_1[24]), .A (n_61), .B (n_50));
AOI21_X1 i_67 (.ZN (n_43), .A (n_317), .B1 (p_0[23]), .B2 (aux[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_261), .B1 (p_0[20]), .B2 (aux[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_318), .B1 (n_261), .B2 (n_63));
OAI21_X1 i_64 (.ZN (n_40), .A (n_314), .B1 (n_259), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_315), .A2 (n_259));
OAI21_X1 i_61 (.ZN (n_37), .A (n_312), .B1 (n_257), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (p_1[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_313), .A2 (n_257));
XOR2_X1 i_58 (.Z (p_1[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (p_1[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (p_1[20]), .A (n_63), .B (n_42));
AOI21_X1 i_55 (.ZN (n_35), .A (n_289), .B1 (p_0[19]), .B2 (aux[19]));
OAI21_X1 i_54 (.ZN (n_34), .A (n_279), .B1 (p_0[16]), .B2 (aux[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_282), .B1 (n_319), .B2 (n_279));
OAI21_X1 i_52 (.ZN (n_32), .A (n_286), .B1 (n_277), .B2 (n_33));
INV_X1 i_51 (.ZN (n_31), .A (n_32));
NOR2_X1 i_50 (.ZN (n_30), .A1 (n_287), .A2 (n_277));
OAI21_X1 i_49 (.ZN (n_29), .A (n_284), .B1 (n_275), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (p_1[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_285), .A2 (n_275));
XOR2_X1 i_46 (.Z (p_1[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (p_1[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (p_1[16]), .A (n_319), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_332), .A2 (n_323));
OAI21_X1 i_42 (.ZN (n_26), .A (n_326), .B1 (p_0[12]), .B2 (aux[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_328), .B1 (n_333), .B2 (n_326));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_331), .B1 (n_325), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_331), .B1 (p_0[13]), .B2 (aux[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (aux[14]), .B1 (n_321), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (p_1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_330), .A2 (n_321));
XOR2_X1 i_34 (.Z (p_1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (p_1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (p_1[12]), .A (n_333), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_346), .A2 (n_337));
AOI21_X1 i_30 (.ZN (n_18), .A (n_342), .B1 (p_0[8]), .B2 (aux[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_342), .B1 (n_347), .B2 (n_340));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_345), .B1 (n_339), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_345), .B1 (p_0[9]), .B2 (aux[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (aux[10]), .B1 (n_335), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (p_1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_344), .A2 (n_335));
XOR2_X1 i_22 (.Z (p_1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (p_1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (p_1[8]), .A (n_347), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_360), .A2 (n_351));
OAI21_X1 i_18 (.ZN (n_10), .A (n_354), .B1 (p_0[4]), .B2 (aux[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_356), .B1 (n_361), .B2 (n_354));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_359), .B1 (n_353), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_359), .B1 (p_0[5]), .B2 (aux[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (aux[6]), .B1 (n_349), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (p_1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_358), .A2 (n_349));
XOR2_X1 i_10 (.Z (p_1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (p_1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (p_1[4]), .A (n_361), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_370), .B1 (n_376), .B2 (n_372));
XOR2_X1 i_6 (.Z (p_1[3]), .A (n_363), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_369), .B1 (p_0[2]), .B2 (aux[2]));
XNOR2_X1 i_4 (.ZN (p_1[2]), .A (n_364), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_365), .B1 (p_0[1]), .B2 (aux[1]));
XOR2_X1 i_2 (.Z (p_1[1]), .A (n_366), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_366), .B1 (p_0[0]), .B2 (aux[0]));
INV_X1 i_0 (.ZN (p_1[0]), .A (n_0));

endmodule //datapath__0_74

module datapath (firstInputComplement, a);

output [31:0] firstInputComplement;
input [31:0] a;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (a[25]));
INV_X1 i_63 (.ZN (n_32), .A (a[21]));
INV_X1 i_62 (.ZN (n_31), .A (a[14]));
INV_X1 i_61 (.ZN (n_30), .A (a[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (a[2]), .A2 (a[1]), .A3 (a[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (a[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (a[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (a[5]), .A3 (a[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (a[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (a[8]), .A3 (a[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (a[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (a[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (a[12]), .A3 (a[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (a[15]), .A3 (a[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (a[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (a[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (a[18]), .A3 (a[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (a[18]), .A3 (a[19]), .A4 (a[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (a[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (a[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (a[23]), .A3 (a[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (a[26]), .A3 (a[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (a[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (a[28]), .A3 (a[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (a[28]), .A3 (a[29]), .A4 (a[30]));
XNOR2_X1 i_35 (.ZN (firstInputComplement[31]), .A (a[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (firstInputComplement[30]), .A (a[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (firstInputComplement[29]), .A (a[29]), .B (n_7));
XOR2_X1 i_32 (.Z (firstInputComplement[28]), .A (a[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (a[27]), .B1 (n_9), .B2 (a[26]));
AND2_X1 i_30 (.ZN (firstInputComplement[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (firstInputComplement[26]), .A (a[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (firstInputComplement[25]), .A (a[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (firstInputComplement[24]), .A (a[24]), .B (n_11));
XOR2_X1 i_26 (.Z (firstInputComplement[23]), .A (a[23]), .B (n_12));
XOR2_X1 i_25 (.Z (firstInputComplement[22]), .A (a[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (firstInputComplement[21]), .A (a[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (firstInputComplement[20]), .A (a[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (firstInputComplement[19]), .A (a[19]), .B (n_16));
XOR2_X1 i_21 (.Z (firstInputComplement[18]), .A (a[18]), .B (n_17));
XOR2_X1 i_20 (.Z (firstInputComplement[17]), .A (a[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (a[16]), .B1 (n_19), .B2 (a[15]));
AND2_X1 i_18 (.ZN (firstInputComplement[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (firstInputComplement[15]), .A (a[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (firstInputComplement[14]), .A (a[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (firstInputComplement[13]), .A (a[13]), .B (n_21));
XOR2_X1 i_14 (.Z (firstInputComplement[12]), .A (a[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (firstInputComplement[11]), .A (a[11]), .B (n_23));
XOR2_X1 i_12 (.Z (firstInputComplement[10]), .A (a[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (a[9]), .B1 (n_25), .B2 (a[8]));
AND2_X1 i_10 (.ZN (firstInputComplement[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (firstInputComplement[8]), .A (a[8]), .B (n_25));
XOR2_X1 i_8 (.Z (firstInputComplement[7]), .A (a[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (a[6]), .B1 (n_27), .B2 (a[5]));
AND2_X1 i_6 (.ZN (firstInputComplement[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (firstInputComplement[5]), .A (a[5]), .B (n_27));
XOR2_X1 i_4 (.Z (firstInputComplement[4]), .A (a[4]), .B (n_28));
XOR2_X1 i_3 (.Z (firstInputComplement[3]), .A (a[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (a[2]), .B1 (a[1]), .B2 (a[0]));
AND2_X1 i_1 (.ZN (firstInputComplement[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (firstInputComplement[1]), .A (a[1]), .B (a[0]));

endmodule //datapath

module radix4Booth (clk_CTS_0_PP_8, clk_CTS_0_PP_14, a, b, clk, reset, en, result, 
    enableOutput);

output enableOutput;
output [63:0] result;
output clk_CTS_0_PP_8;
input [31:0] a;
input [31:0] b;
input clk;
input en;
input reset;
input clk_CTS_0_PP_14;
wire CTS_n_tid0_189;
wire \firstInputComplement[31] ;
wire \firstInputComplement[30] ;
wire \firstInputComplement[29] ;
wire \firstInputComplement[28] ;
wire \firstInputComplement[27] ;
wire \firstInputComplement[26] ;
wire \firstInputComplement[25] ;
wire \firstInputComplement[24] ;
wire \firstInputComplement[23] ;
wire \firstInputComplement[22] ;
wire \firstInputComplement[21] ;
wire \firstInputComplement[20] ;
wire \firstInputComplement[19] ;
wire \firstInputComplement[18] ;
wire \firstInputComplement[17] ;
wire \firstInputComplement[16] ;
wire \firstInputComplement[15] ;
wire \firstInputComplement[14] ;
wire \firstInputComplement[13] ;
wire \firstInputComplement[12] ;
wire \firstInputComplement[11] ;
wire \firstInputComplement[10] ;
wire \firstInputComplement[9] ;
wire \firstInputComplement[8] ;
wire \firstInputComplement[7] ;
wire \firstInputComplement[6] ;
wire \firstInputComplement[5] ;
wire \firstInputComplement[4] ;
wire \firstInputComplement[3] ;
wire \firstInputComplement[2] ;
wire \firstInputComplement[1] ;
wire hfn_ipo_n17;
wire n_1_3;
wire n_1_0;
wire n_1_4;
wire n_1_1;
wire n_1_5;
wire n_1_2;
wire n_1_6;
wire n_1_7;
wire n_1_8;
wire n_1_9;
wire n_1_10;
wire n_1_11;
wire n_1_12;
wire n_1_13;
wire n_1_14;
wire n_1_15;
wire n_1_16;
wire n_1_17;
wire n_1_18;
wire n_1_19;
wire n_1_20;
wire n_1_21;
wire n_1_22;
wire n_1_23;
wire n_1_24;
wire n_1_25;
wire n_1_26;
wire n_1_27;
wire n_1_28;
wire n_1_29;
wire n_1_30;
wire n_1_31;
wire n_1_32;
wire n_1_33;
wire n_1_34;
wire n_1_35;
wire n_1_36;
wire n_1_37;
wire n_1_38;
wire n_1_39;
wire n_1_40;
wire n_1_41;
wire n_1_42;
wire n_1_43;
wire n_1_44;
wire n_1_45;
wire n_1_46;
wire n_1_47;
wire n_1_48;
wire n_1_49;
wire n_1_50;
wire n_1_51;
wire n_1_52;
wire n_1_53;
wire n_1_54;
wire n_1_55;
wire n_1_56;
wire n_1_57;
wire n_1_58;
wire n_1_59;
wire n_1_60;
wire n_1_61;
wire n_1_62;
wire n_1_63;
wire n_1_64;
wire n_1_65;
wire n_1_66;
wire n_1_67;
wire n_1_68;
wire n_1_69;
wire n_1_70;
wire n_1_71;
wire n_1_72;
wire n_1_73;
wire n_1_74;
wire n_1_75;
wire n_1_76;
wire n_1_77;
wire n_1_78;
wire n_1_79;
wire n_1_80;
wire n_1_81;
wire n_1_82;
wire n_1_83;
wire n_1_84;
wire n_1_85;
wire n_1_86;
wire n_1_87;
wire n_1_88;
wire n_1_89;
wire n_1_90;
wire n_1_91;
wire n_1_92;
wire n_1_93;
wire n_1_94;
wire n_1_95;
wire n_1_96;
wire n_1_97;
wire n_1_98;
wire n_1_99;
wire n_1_100;
wire n_1_101;
wire n_1_102;
wire n_1_103;
wire n_1_104;
wire n_1_105;
wire n_1_106;
wire n_1_107;
wire n_1_108;
wire n_1_109;
wire n_1_110;
wire n_1_111;
wire n_1_112;
wire n_1_113;
wire n_1_114;
wire n_1_115;
wire n_1_116;
wire n_1_117;
wire n_1_118;
wire n_1_119;
wire n_1_120;
wire n_1_121;
wire n_1_122;
wire n_1_123;
wire n_1_124;
wire n_1_125;
wire n_1_126;
wire n_1_127;
wire n_1_128;
wire n_1_129;
wire n_1_130;
wire n_1_131;
wire n_1_132;
wire n_1_133;
wire n_1_134;
wire n_1_135;
wire n_1_136;
wire n_1_137;
wire n_1_138;
wire n_1_139;
wire n_1_140;
wire n_1_141;
wire n_1_142;
wire n_1_143;
wire n_1_144;
wire n_1_145;
wire n_1_146;
wire n_1_147;
wire n_1_148;
wire n_1_149;
wire n_1_150;
wire n_1_151;
wire n_1_152;
wire n_1_153;
wire n_1_154;
wire n_1_155;
wire n_1_156;
wire n_1_157;
wire n_1_158;
wire n_1_159;
wire n_1_160;
wire n_1_161;
wire n_1_162;
wire n_1_163;
wire n_1_164;
wire n_1_165;
wire n_1_166;
wire n_1_167;
wire n_1_168;
wire n_1_169;
wire n_1_170;
wire n_1_171;
wire n_1_172;
wire n_1_173;
wire n_1_174;
wire n_1_175;
wire n_1_176;
wire n_1_177;
wire n_1_178;
wire n_1_179;
wire n_1_180;
wire n_1_181;
wire n_1_182;
wire n_1_183;
wire n_1_184;
wire n_1_185;
wire n_1_186;
wire n_1_187;
wire n_1_188;
wire n_1_189;
wire n_1_190;
wire n_1_191;
wire n_1_192;
wire n_1_193;
wire n_1_194;
wire n_1_195;
wire n_1_196;
wire n_1_197;
wire n_1_198;
wire n_1_199;
wire n_1_200;
wire n_1_201;
wire n_1_202;
wire n_1_203;
wire n_1_204;
wire n_1_205;
wire n_1_206;
wire n_1_207;
wire n_1_208;
wire n_1_209;
wire n_1_210;
wire n_1_211;
wire n_1_212;
wire n_1_213;
wire n_1_214;
wire n_1_215;
wire n_1_216;
wire n_1_217;
wire n_1_218;
wire n_1_219;
wire n_1_220;
wire n_1_221;
wire n_1_222;
wire n_1_223;
wire n_1_224;
wire n_1_225;
wire n_1_226;
wire n_1_227;
wire n_1_228;
wire n_1_229;
wire n_1_230;
wire n_1_231;
wire n_1_232;
wire n_1_233;
wire n_1_234;
wire n_1_235;
wire n_1_236;
wire n_1_237;
wire n_1_238;
wire n_1_239;
wire n_1_240;
wire n_1_241;
wire n_1_242;
wire n_1_243;
wire n_1_244;
wire n_1_245;
wire n_1_246;
wire n_1_247;
wire n_1_248;
wire n_1_249;
wire n_1_250;
wire n_1_251;
wire n_1_252;
wire n_1_253;
wire n_1_254;
wire n_1_255;
wire n_1_256;
wire n_1_257;
wire n_1_258;
wire n_1_259;
wire n_1_260;
wire n_1_261;
wire n_1_262;
wire n_1_263;
wire n_1_264;
wire n_1_265;
wire n_1_266;
wire n_1_267;
wire n_1_268;
wire n_1_269;
wire n_1_270;
wire n_1_271;
wire n_1_272;
wire n_1_273;
wire n_1_274;
wire n_1_275;
wire n_1_276;
wire n_1_277;
wire n_1_278;
wire n_1_279;
wire n_1_280;
wire n_1_281;
wire n_1_282;
wire n_1_283;
wire n_1_284;
wire n_1_285;
wire n_1_286;
wire n_1_287;
wire n_1_288;
wire n_1_289;
wire n_1_290;
wire n_1_291;
wire n_1_292;
wire n_1_293;
wire n_1_294;
wire n_1_295;
wire n_1_296;
wire n_1_297;
wire n_1_298;
wire n_1_299;
wire n_1_300;
wire n_1_301;
wire n_1_302;
wire n_1_303;
wire n_1_304;
wire n_1_305;
wire n_1_306;
wire n_1_307;
wire n_1_308;
wire n_1_309;
wire n_1_310;
wire n_1_311;
wire n_1_312;
wire n_1_313;
wire n_1_314;
wire n_1_315;
wire n_1_316;
wire n_1_317;
wire n_1_318;
wire n_1_319;
wire n_1_320;
wire n_1_321;
wire n_1_322;
wire n_1_323;
wire n_1_324;
wire n_1_325;
wire n_1_326;
wire n_1_327;
wire n_1_328;
wire n_1_329;
wire n_1_330;
wire n_1_331;
wire n_1_332;
wire n_1_333;
wire n_1_334;
wire n_1_335;
wire n_1_336;
wire n_1_337;
wire n_1_338;
wire n_1_339;
wire n_1_340;
wire n_1_341;
wire n_1_342;
wire n_1_343;
wire n_1_344;
wire n_1_345;
wire n_1_346;
wire n_1_347;
wire n_1_348;
wire n_1_349;
wire n_1_350;
wire n_1_351;
wire n_1_352;
wire n_1_353;
wire n_1_354;
wire n_1_355;
wire n_1_356;
wire n_1_357;
wire n_1_358;
wire n_1_359;
wire n_1_360;
wire n_1_361;
wire n_1_362;
wire n_1_363;
wire n_1_364;
wire n_1_365;
wire n_1_366;
wire n_1_367;
wire n_1_368;
wire n_1_369;
wire n_1_370;
wire n_1_371;
wire n_1_372;
wire n_1_373;
wire n_1_374;
wire n_1_375;
wire n_1_376;
wire n_1_377;
wire n_1_378;
wire n_1_379;
wire n_1_380;
wire n_1_381;
wire n_1_382;
wire n_1_383;
wire n_1_384;
wire n_1_385;
wire n_1_386;
wire n_1_387;
wire n_1_388;
wire n_1_389;
wire n_1_390;
wire n_1_391;
wire n_1_392;
wire n_1_393;
wire n_1_394;
wire n_1_395;
wire n_1_396;
wire n_1_397;
wire n_1_398;
wire n_1_399;
wire n_1_400;
wire n_1_401;
wire n_1_402;
wire n_1_403;
wire n_1_404;
wire n_1_405;
wire n_1_406;
wire n_1_407;
wire n_1_408;
wire n_1_409;
wire n_1_410;
wire n_1_411;
wire n_1_412;
wire n_1_413;
wire n_1_414;
wire n_1_415;
wire n_1_416;
wire n_1_417;
wire n_1_418;
wire n_1_419;
wire n_1_420;
wire n_1_421;
wire n_1_422;
wire n_1_423;
wire n_1_424;
wire n_1_425;
wire n_1_426;
wire n_1_427;
wire n_1_428;
wire n_1_429;
wire n_1_430;
wire n_1_431;
wire n_1_432;
wire n_1_433;
wire n_1_434;
wire n_1_435;
wire n_1_436;
wire n_1_437;
wire n_1_438;
wire n_1_439;
wire n_1_440;
wire n_1_441;
wire n_1_442;
wire n_1_443;
wire n_1_444;
wire n_1_445;
wire n_1_446;
wire n_1_447;
wire n_1_448;
wire n_1_449;
wire n_1_450;
wire n_1_451;
wire n_1_452;
wire n_1_453;
wire n_1_454;
wire n_1_455;
wire n_1_456;
wire n_1_457;
wire n_1_458;
wire n_1_459;
wire n_1_460;
wire n_1_461;
wire n_1_462;
wire n_1_463;
wire n_1_464;
wire n_1_465;
wire n_1_466;
wire n_1_467;
wire n_1_468;
wire n_1_469;
wire n_1_470;
wire n_1_471;
wire n_1_472;
wire n_1_473;
wire n_1_474;
wire n_1_475;
wire n_1_476;
wire n_1_477;
wire n_1_478;
wire n_1_479;
wire n_1_480;
wire n_1_481;
wire n_1_482;
wire n_1_483;
wire n_1_484;
wire n_1_485;
wire n_1_486;
wire n_1_487;
wire n_1_488;
wire n_1_489;
wire n_1_490;
wire n_1_491;
wire n_1_492;
wire n_1_493;
wire n_1_494;
wire n_1_495;
wire n_1_496;
wire n_1_497;
wire n_1_498;
wire n_1_499;
wire n_1_500;
wire n_1_501;
wire n_1_502;
wire n_1_503;
wire n_1_504;
wire n_1_505;
wire n_1_506;
wire n_1_507;
wire n_1_508;
wire n_1_509;
wire n_1_510;
wire n_1_511;
wire n_1_512;
wire n_1_513;
wire n_1_514;
wire n_1_515;
wire n_1_516;
wire n_1_517;
wire n_1_518;
wire n_1_519;
wire n_1_520;
wire n_1_521;
wire n_1_522;
wire n_1_523;
wire n_1_524;
wire n_1_525;
wire n_1_526;
wire n_1_527;
wire n_1_528;
wire n_1_529;
wire n_1_530;
wire n_1_531;
wire n_1_532;
wire n_1_533;
wire n_1_534;
wire n_1_535;
wire n_1_536;
wire n_1_537;
wire n_1_538;
wire n_1_539;
wire n_1_540;
wire n_1_541;
wire n_1_542;
wire n_1_543;
wire n_1_544;
wire n_1_545;
wire n_1_546;
wire n_1_547;
wire n_1_548;
wire n_1_549;
wire n_1_550;
wire n_1_551;
wire n_1_552;
wire n_1_553;
wire n_1_554;
wire n_1_555;
wire n_1_556;
wire n_1_557;
wire n_1_558;
wire n_1_559;
wire n_1_560;
wire n_1_561;
wire n_1_562;
wire n_1_563;
wire n_1_564;
wire n_1_565;
wire n_1_566;
wire n_1_567;
wire n_1_568;
wire n_1_569;
wire n_1_570;
wire n_1_571;
wire n_1_572;
wire n_1_573;
wire n_1_574;
wire n_1_575;
wire n_1_576;
wire n_1_577;
wire n_1_578;
wire n_1_579;
wire n_1_580;
wire n_1_581;
wire n_1_582;
wire n_1_583;
wire n_1_584;
wire n_1_585;
wire n_1_586;
wire n_1_587;
wire n_1_588;
wire n_1_589;
wire n_1_590;
wire n_1_591;
wire n_1_592;
wire n_1_593;
wire n_1_594;
wire n_1_595;
wire n_1_596;
wire n_1_597;
wire n_1_598;
wire n_1_599;
wire n_1_600;
wire n_1_601;
wire n_1_602;
wire n_1_603;
wire n_1_604;
wire n_1_605;
wire n_1_606;
wire n_1_607;
wire n_1_608;
wire n_1_609;
wire n_1_610;
wire n_1_611;
wire n_1_612;
wire n_1_613;
wire n_1_614;
wire n_1_615;
wire n_1_616;
wire n_1_617;
wire n_1_618;
wire n_1_619;
wire n_1_620;
wire n_1_621;
wire n_1_622;
wire n_1_623;
wire n_1_624;
wire n_1_625;
wire n_1_626;
wire n_1_627;
wire n_1_628;
wire n_1_629;
wire n_1_630;
wire n_1_631;
wire n_1_632;
wire n_1_633;
wire n_1_634;
wire n_1_635;
wire n_1_636;
wire n_1_637;
wire n_1_638;
wire n_1_639;
wire n_1_640;
wire n_1_641;
wire n_1_642;
wire n_1_643;
wire n_1_644;
wire n_1_645;
wire n_1_646;
wire n_1_647;
wire n_1_648;
wire n_1_649;
wire n_1_650;
wire n_1_651;
wire n_1_652;
wire n_1_653;
wire n_1_654;
wire n_1_655;
wire n_1_656;
wire n_1_657;
wire n_1_658;
wire n_1_659;
wire n_1_660;
wire n_1_661;
wire n_1_662;
wire n_1_663;
wire n_1_664;
wire n_1_665;
wire n_1_666;
wire n_1_667;
wire n_1_668;
wire n_1_669;
wire n_1_670;
wire n_1_671;
wire n_1_672;
wire n_1_673;
wire n_1_674;
wire n_1_675;
wire n_1_676;
wire n_1_677;
wire n_1_678;
wire n_1_679;
wire n_1_680;
wire n_1_681;
wire n_1_682;
wire n_1_683;
wire n_1_684;
wire n_1_685;
wire n_1_686;
wire n_1_687;
wire n_1_688;
wire n_1_689;
wire n_1_690;
wire n_1_691;
wire n_1_692;
wire n_1_693;
wire n_1_694;
wire n_1_695;
wire n_1_696;
wire n_1_697;
wire n_1_698;
wire n_1_699;
wire n_1_700;
wire n_1_701;
wire n_1_702;
wire n_1_703;
wire n_1_704;
wire n_1_705;
wire n_1_706;
wire n_1_707;
wire n_1_708;
wire n_1_709;
wire n_1_710;
wire n_1_711;
wire n_1_712;
wire n_1_713;
wire n_1_714;
wire n_1_715;
wire n_1_716;
wire n_1_717;
wire n_1_718;
wire n_1_719;
wire n_1_720;
wire n_1_721;
wire n_1_722;
wire n_1_723;
wire n_1_724;
wire n_1_725;
wire n_1_726;
wire n_1_727;
wire n_1_728;
wire n_1_729;
wire n_1_730;
wire n_1_731;
wire n_1_732;
wire n_1_733;
wire n_1_734;
wire n_1_735;
wire n_1_736;
wire n_1_737;
wire n_1_738;
wire n_1_739;
wire n_1_740;
wire n_1_741;
wire n_1_742;
wire n_1_743;
wire n_1_744;
wire n_1_745;
wire n_1_746;
wire n_1_747;
wire n_1_748;
wire n_1_749;
wire n_1_750;
wire n_1_751;
wire n_1_752;
wire n_1_753;
wire n_1_754;
wire n_1_755;
wire n_1_756;
wire n_1_757;
wire n_1_758;
wire n_1_759;
wire n_1_760;
wire n_1_761;
wire n_1_762;
wire n_1_763;
wire n_1_764;
wire n_1_765;
wire n_1_766;
wire n_1_767;
wire n_1_768;
wire n_1_769;
wire n_1_770;
wire n_1_771;
wire n_1_772;
wire n_1_773;
wire n_1_774;
wire n_1_775;
wire n_1_776;
wire n_1_777;
wire n_1_778;
wire n_1_779;
wire n_1_780;
wire n_1_781;
wire n_1_782;
wire n_1_783;
wire n_1_784;
wire n_1_785;
wire n_1_786;
wire n_1_787;
wire n_1_788;
wire n_1_789;
wire n_1_790;
wire n_1_791;
wire n_1_792;
wire n_1_793;
wire n_1_794;
wire n_1_795;
wire n_1_796;
wire n_1_797;
wire n_1_798;
wire n_1_799;
wire n_1_800;
wire n_1_801;
wire n_1_802;
wire n_1_803;
wire n_1_804;
wire n_1_805;
wire n_1_806;
wire n_1_807;
wire n_1_808;
wire n_1_809;
wire n_1_810;
wire n_1_811;
wire n_1_812;
wire n_1_813;
wire n_1_814;
wire n_1_815;
wire n_1_816;
wire n_1_817;
wire n_1_818;
wire n_1_819;
wire n_1_820;
wire n_1_821;
wire n_1_822;
wire n_1_823;
wire n_1_824;
wire n_1_825;
wire n_1_826;
wire n_1_827;
wire n_1_828;
wire n_1_829;
wire n_1_830;
wire n_1_831;
wire n_1_832;
wire n_1_833;
wire n_1_834;
wire n_1_835;
wire n_1_836;
wire n_1_837;
wire n_1_838;
wire n_1_839;
wire n_1_840;
wire n_1_841;
wire n_1_842;
wire n_1_843;
wire n_1_844;
wire n_1_845;
wire n_1_846;
wire n_1_847;
wire n_1_848;
wire n_1_849;
wire n_1_850;
wire n_1_851;
wire n_1_852;
wire n_1_853;
wire n_1_854;
wire n_1_855;
wire n_1_856;
wire n_1_857;
wire n_1_858;
wire n_1_859;
wire n_1_860;
wire n_1_861;
wire n_1_862;
wire n_1_863;
wire n_1_864;
wire n_1_865;
wire n_1_866;
wire n_1_867;
wire n_1_868;
wire n_1_869;
wire n_1_870;
wire n_1_871;
wire n_1_872;
wire n_1_873;
wire n_1_874;
wire n_1_875;
wire n_1_876;
wire n_1_877;
wire n_1_878;
wire n_1_879;
wire n_1_880;
wire n_1_881;
wire n_1_882;
wire n_1_883;
wire n_1_884;
wire n_1_885;
wire n_1_886;
wire n_1_887;
wire n_1_888;
wire n_1_889;
wire n_1_890;
wire n_1_891;
wire n_1_892;
wire n_1_893;
wire n_1_894;
wire n_1_895;
wire n_1_896;
wire n_1_897;
wire n_1_898;
wire n_1_899;
wire n_1_900;
wire n_1_901;
wire n_1_902;
wire n_1_903;
wire n_1_904;
wire n_1_905;
wire n_1_906;
wire n_1_907;
wire n_1_908;
wire n_1_909;
wire n_1_910;
wire n_1_911;
wire n_1_912;
wire n_1_913;
wire n_1_914;
wire n_1_915;
wire n_1_916;
wire n_1_917;
wire n_1_918;
wire n_1_919;
wire n_1_920;
wire n_1_921;
wire n_1_922;
wire n_1_923;
wire n_1_924;
wire n_1_925;
wire n_1_926;
wire n_1_927;
wire n_1_928;
wire n_1_929;
wire n_1_930;
wire n_1_931;
wire n_1_932;
wire n_1_933;
wire n_1_934;
wire n_1_935;
wire n_1_936;
wire n_1_937;
wire n_1_938;
wire \counter[4] ;
wire \counter[3] ;
wire \counter[2] ;
wire \counter[1] ;
wire \counter[0] ;
wire resetReg;
wire \aux[63] ;
wire \aux[62] ;
wire \aux[61] ;
wire \aux[60] ;
wire \aux[59] ;
wire \aux[58] ;
wire \aux[57] ;
wire \aux[56] ;
wire \aux[55] ;
wire \aux[54] ;
wire \aux[53] ;
wire \aux[52] ;
wire \aux[51] ;
wire \aux[50] ;
wire \aux[49] ;
wire \aux[48] ;
wire \aux[47] ;
wire \aux[46] ;
wire \aux[45] ;
wire \aux[44] ;
wire \aux[43] ;
wire \aux[42] ;
wire \aux[41] ;
wire \aux[40] ;
wire \aux[39] ;
wire \aux[38] ;
wire \aux[37] ;
wire \aux[36] ;
wire \aux[35] ;
wire \aux[34] ;
wire \aux[33] ;
wire \aux[32] ;
wire \aux[31] ;
wire \aux[30] ;
wire \aux[29] ;
wire \aux[28] ;
wire \aux[27] ;
wire \aux[26] ;
wire \aux[25] ;
wire \aux[24] ;
wire \aux[23] ;
wire \aux[22] ;
wire \aux[21] ;
wire \aux[20] ;
wire \aux[19] ;
wire \aux[18] ;
wire \aux[17] ;
wire \aux[16] ;
wire \aux[15] ;
wire \aux[14] ;
wire \aux[13] ;
wire \aux[12] ;
wire \aux[11] ;
wire \aux[10] ;
wire \aux[9] ;
wire \aux[8] ;
wire \aux[7] ;
wire \aux[6] ;
wire \aux[5] ;
wire \aux[4] ;
wire \aux[3] ;
wire \aux[2] ;
wire \aux[1] ;
wire \aux[0] ;
wire uc_0;
wire n_268;
wire n_264;
wire n_263;
wire n_262;
wire n_261;
wire n_260;
wire n_259;
wire n_258;
wire n_257;
wire n_256;
wire n_255;
wire n_254;
wire n_253;
wire n_252;
wire n_251;
wire n_250;
wire n_249;
wire n_248;
wire n_247;
wire n_246;
wire n_245;
wire n_244;
wire n_243;
wire n_242;
wire n_241;
wire n_240;
wire n_239;
wire n_238;
wire n_237;
wire n_236;
wire n_235;
wire n_234;
wire n_233;
wire n_232;
wire n_231;
wire n_230;
wire n_229;
wire n_228;
wire n_227;
wire n_226;
wire n_225;
wire n_224;
wire n_223;
wire n_222;
wire n_221;
wire n_220;
wire n_219;
wire n_218;
wire n_217;
wire n_216;
wire n_215;
wire n_214;
wire n_213;
wire n_212;
wire n_211;
wire n_210;
wire n_209;
wire n_208;
wire n_207;
wire n_206;
wire n_205;
wire n_204;
wire n_203;
wire n_202;
wire n_201;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_67;
wire n_267;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_265;
wire n_266;
wire CTS_n_tid0_81;
wire n_1;
wire n_269;
wire CTS_n_tid0_84;
wire CTS_n_tid0_82;
wire hfn_ipo_n15;
wire hfn_ipo_n16;
wire hfn_ipo_n13;
wire hfn_ipo_n14;
wire drc_ipo_n19;
wire CTS_n_tid0_153;
wire CTS_n_tid1_73;
wire CLOCK_sgo__n273;
wire CTS_n_tid1_76;
wire CTS_n_tid0_247;
wire CTS_n_tid0_206;


DFF_X1 \aux_reg[0]  (.Q (\aux[0] ), .CK (CTS_n_tid1_76), .D (n_137));
DFF_X1 \aux_reg[1]  (.Q (\aux[1] ), .CK (CTS_n_tid1_76), .D (n_138));
DFF_X1 \aux_reg[2]  (.Q (\aux[2] ), .CK (CTS_n_tid1_76), .D (n_139));
DFF_X1 \aux_reg[3]  (.Q (\aux[3] ), .CK (CTS_n_tid1_76), .D (n_140));
DFF_X1 \aux_reg[4]  (.Q (\aux[4] ), .CK (CTS_n_tid1_76), .D (n_141));
DFF_X1 \aux_reg[5]  (.Q (\aux[5] ), .CK (CTS_n_tid1_76), .D (n_142));
DFF_X1 \aux_reg[6]  (.Q (\aux[6] ), .CK (CTS_n_tid1_76), .D (n_143));
DFF_X1 \aux_reg[7]  (.Q (\aux[7] ), .CK (CTS_n_tid1_76), .D (n_144));
DFF_X1 \aux_reg[8]  (.Q (\aux[8] ), .CK (CTS_n_tid1_76), .D (n_145));
DFF_X1 \aux_reg[9]  (.Q (\aux[9] ), .CK (CTS_n_tid1_76), .D (n_146));
DFF_X1 \aux_reg[10]  (.Q (\aux[10] ), .CK (CTS_n_tid1_76), .D (n_147));
DFF_X1 \aux_reg[11]  (.Q (\aux[11] ), .CK (CTS_n_tid1_76), .D (n_148));
DFF_X1 \aux_reg[12]  (.Q (\aux[12] ), .CK (CTS_n_tid1_76), .D (n_149));
DFF_X1 \aux_reg[13]  (.Q (\aux[13] ), .CK (CTS_n_tid1_76), .D (n_150));
DFF_X1 \aux_reg[14]  (.Q (\aux[14] ), .CK (CTS_n_tid1_76), .D (n_151));
DFF_X1 \aux_reg[15]  (.Q (\aux[15] ), .CK (CTS_n_tid1_76), .D (n_152));
DFF_X1 \aux_reg[16]  (.Q (\aux[16] ), .CK (CTS_n_tid1_76), .D (n_153));
DFF_X1 \aux_reg[17]  (.Q (\aux[17] ), .CK (CTS_n_tid1_76), .D (n_154));
DFF_X1 \aux_reg[18]  (.Q (\aux[18] ), .CK (CTS_n_tid1_76), .D (n_155));
DFF_X1 \aux_reg[19]  (.Q (\aux[19] ), .CK (CTS_n_tid1_76), .D (n_156));
DFF_X1 \aux_reg[20]  (.Q (\aux[20] ), .CK (CTS_n_tid1_76), .D (n_157));
DFF_X1 \aux_reg[21]  (.Q (\aux[21] ), .CK (CTS_n_tid1_76), .D (n_158));
DFF_X1 \aux_reg[22]  (.Q (\aux[22] ), .CK (CTS_n_tid1_76), .D (n_159));
DFF_X1 \aux_reg[23]  (.Q (\aux[23] ), .CK (CTS_n_tid1_76), .D (n_160));
DFF_X1 \aux_reg[24]  (.Q (\aux[24] ), .CK (CTS_n_tid1_76), .D (n_161));
DFF_X1 \aux_reg[25]  (.Q (\aux[25] ), .CK (CTS_n_tid1_76), .D (n_162));
DFF_X1 \aux_reg[26]  (.Q (\aux[26] ), .CK (CTS_n_tid1_76), .D (n_163));
DFF_X1 \aux_reg[27]  (.Q (\aux[27] ), .CK (CTS_n_tid1_76), .D (n_164));
DFF_X1 \aux_reg[28]  (.Q (\aux[28] ), .CK (CTS_n_tid1_76), .D (n_165));
DFF_X1 \aux_reg[29]  (.Q (\aux[29] ), .CK (CTS_n_tid1_76), .D (n_166));
DFF_X1 \aux_reg[30]  (.Q (\aux[30] ), .CK (CTS_n_tid1_76), .D (n_167));
DFF_X1 \aux_reg[31]  (.Q (\aux[31] ), .CK (CTS_n_tid1_76), .D (n_168));
DFF_X1 \aux_reg[32]  (.Q (\aux[32] ), .CK (CTS_n_tid1_76), .D (n_169));
DFF_X1 \aux_reg[33]  (.Q (\aux[33] ), .CK (CTS_n_tid1_76), .D (n_170));
DFF_X1 \aux_reg[34]  (.Q (\aux[34] ), .CK (CTS_n_tid1_76), .D (n_171));
DFF_X1 \aux_reg[35]  (.Q (\aux[35] ), .CK (CTS_n_tid1_76), .D (n_172));
DFF_X1 \aux_reg[36]  (.Q (\aux[36] ), .CK (CTS_n_tid1_76), .D (n_173));
DFF_X1 \aux_reg[37]  (.Q (\aux[37] ), .CK (CTS_n_tid1_76), .D (n_174));
DFF_X1 \aux_reg[38]  (.Q (\aux[38] ), .CK (CTS_n_tid1_76), .D (n_175));
DFF_X1 \aux_reg[39]  (.Q (\aux[39] ), .CK (CTS_n_tid1_76), .D (n_176));
DFF_X1 \aux_reg[40]  (.Q (\aux[40] ), .CK (CTS_n_tid1_76), .D (n_177));
DFF_X1 \aux_reg[41]  (.Q (\aux[41] ), .CK (CTS_n_tid1_76), .D (n_178));
DFF_X1 \aux_reg[42]  (.Q (\aux[42] ), .CK (CTS_n_tid1_76), .D (n_179));
DFF_X1 \aux_reg[43]  (.Q (\aux[43] ), .CK (CTS_n_tid1_76), .D (n_180));
DFF_X1 \aux_reg[44]  (.Q (\aux[44] ), .CK (CTS_n_tid1_76), .D (n_181));
DFF_X1 \aux_reg[45]  (.Q (\aux[45] ), .CK (CTS_n_tid1_76), .D (n_182));
DFF_X1 \aux_reg[46]  (.Q (\aux[46] ), .CK (CTS_n_tid1_76), .D (n_183));
DFF_X1 \aux_reg[47]  (.Q (\aux[47] ), .CK (CTS_n_tid1_76), .D (n_184));
DFF_X1 \aux_reg[48]  (.Q (\aux[48] ), .CK (CTS_n_tid1_76), .D (n_185));
DFF_X1 \aux_reg[49]  (.Q (\aux[49] ), .CK (CTS_n_tid1_76), .D (n_186));
DFF_X1 \aux_reg[50]  (.Q (\aux[50] ), .CK (CTS_n_tid1_76), .D (n_187));
DFF_X1 \aux_reg[51]  (.Q (\aux[51] ), .CK (CTS_n_tid1_76), .D (n_188));
DFF_X1 \aux_reg[52]  (.Q (\aux[52] ), .CK (CTS_n_tid1_76), .D (n_189));
DFF_X1 \aux_reg[53]  (.Q (\aux[53] ), .CK (CTS_n_tid1_76), .D (n_190));
DFF_X1 \aux_reg[54]  (.Q (\aux[54] ), .CK (CTS_n_tid1_76), .D (n_191));
DFF_X1 \aux_reg[55]  (.Q (\aux[55] ), .CK (CTS_n_tid1_76), .D (n_192));
DFF_X1 \aux_reg[56]  (.Q (\aux[56] ), .CK (CTS_n_tid1_76), .D (n_193));
DFF_X1 \aux_reg[57]  (.Q (\aux[57] ), .CK (CTS_n_tid1_76), .D (n_194));
DFF_X1 \aux_reg[58]  (.Q (\aux[58] ), .CK (CTS_n_tid1_76), .D (n_195));
DFF_X1 \aux_reg[59]  (.Q (\aux[59] ), .CK (CTS_n_tid1_76), .D (n_196));
DFF_X1 \aux_reg[60]  (.Q (\aux[60] ), .CK (CTS_n_tid1_76), .D (n_197));
DFF_X1 \aux_reg[61]  (.Q (\aux[61] ), .CK (CTS_n_tid1_76), .D (n_198));
DFF_X1 \aux_reg[62]  (.Q (\aux[62] ), .CK (CTS_n_tid1_76), .D (n_199));
DFF_X1 \aux_reg[63]  (.Q (\aux[63] ), .CK (CTS_n_tid1_76), .D (n_200));
CLKGATETST_X4 clk_gate_aux_reg (.GCK (CTS_n_tid1_73), .CK (CTS_n_tid0_189), .E (n_265), .SE (1'b0 ));
MUX2_X1 resetReg_reg_enable_mux_0 (.Z (n_269), .A (resetReg), .B (n_67), .S (n_267));
DFF_X1 resetReg_reg (.Q (resetReg), .CK (CTS_n_tid0_153), .D (n_269));
DFF_X1 \counter_reg[0]  (.Q (\counter[0] ), .CK (n_1), .D (n_132));
DFF_X1 \counter_reg[1]  (.Q (\counter[1] ), .CK (n_1), .D (n_133));
DFF_X1 \counter_reg[2]  (.Q (\counter[2] ), .CK (n_1), .D (n_134));
DFF_X1 \counter_reg[3]  (.Q (\counter[3] ), .CK (n_1), .D (n_135));
DFF_X1 \counter_reg[4]  (.Q (\counter[4] ), .CK (n_1), .D (n_136));
CLKGATETST_X1 clk_gate_counter_reg (.GCK (n_1), .CK (CTS_n_tid0_153), .E (en), .SE (1'b0 ));
DFF_X1 \result_reg[0]  (.Q (result[0]), .CK (CTS_n_tid0_81), .D (n_68));
DFF_X1 \result_reg[1]  (.Q (result[1]), .CK (CTS_n_tid0_81), .D (n_69));
DFF_X1 \result_reg[2]  (.Q (result[2]), .CK (CTS_n_tid0_81), .D (n_70));
DFF_X1 \result_reg[3]  (.Q (result[3]), .CK (CTS_n_tid0_81), .D (n_71));
DFF_X1 \result_reg[4]  (.Q (result[4]), .CK (CTS_n_tid0_81), .D (n_72));
DFF_X1 \result_reg[5]  (.Q (result[5]), .CK (CTS_n_tid0_81), .D (n_73));
DFF_X1 \result_reg[6]  (.Q (result[6]), .CK (CTS_n_tid0_81), .D (n_74));
DFF_X1 \result_reg[7]  (.Q (result[7]), .CK (CTS_n_tid0_81), .D (n_75));
DFF_X1 \result_reg[8]  (.Q (result[8]), .CK (CTS_n_tid0_81), .D (n_76));
DFF_X1 \result_reg[9]  (.Q (result[9]), .CK (CTS_n_tid0_81), .D (n_77));
DFF_X1 \result_reg[10]  (.Q (result[10]), .CK (CTS_n_tid0_81), .D (n_78));
DFF_X1 \result_reg[11]  (.Q (result[11]), .CK (CTS_n_tid0_81), .D (n_79));
DFF_X1 \result_reg[12]  (.Q (result[12]), .CK (CTS_n_tid0_81), .D (n_80));
DFF_X1 \result_reg[13]  (.Q (result[13]), .CK (CTS_n_tid0_81), .D (n_81));
DFF_X1 \result_reg[14]  (.Q (result[14]), .CK (CTS_n_tid0_81), .D (n_82));
DFF_X1 \result_reg[15]  (.Q (result[15]), .CK (CTS_n_tid0_81), .D (n_83));
DFF_X1 \result_reg[16]  (.Q (result[16]), .CK (CTS_n_tid0_81), .D (n_84));
DFF_X1 \result_reg[17]  (.Q (result[17]), .CK (CTS_n_tid0_81), .D (n_85));
DFF_X1 \result_reg[18]  (.Q (result[18]), .CK (CTS_n_tid0_81), .D (n_86));
DFF_X1 \result_reg[19]  (.Q (result[19]), .CK (CTS_n_tid0_81), .D (n_87));
DFF_X1 \result_reg[20]  (.Q (result[20]), .CK (CTS_n_tid0_81), .D (n_88));
DFF_X1 \result_reg[21]  (.Q (result[21]), .CK (CTS_n_tid0_81), .D (n_89));
DFF_X1 \result_reg[22]  (.Q (result[22]), .CK (CTS_n_tid0_81), .D (n_90));
DFF_X1 \result_reg[23]  (.Q (result[23]), .CK (CTS_n_tid0_81), .D (n_91));
DFF_X1 \result_reg[24]  (.Q (result[24]), .CK (CTS_n_tid0_81), .D (n_92));
DFF_X1 \result_reg[25]  (.Q (result[25]), .CK (CTS_n_tid0_81), .D (n_93));
DFF_X1 \result_reg[26]  (.Q (result[26]), .CK (CTS_n_tid0_81), .D (n_94));
DFF_X1 \result_reg[27]  (.Q (result[27]), .CK (CTS_n_tid0_81), .D (n_95));
DFF_X1 \result_reg[28]  (.Q (result[28]), .CK (CTS_n_tid0_81), .D (n_96));
DFF_X1 \result_reg[29]  (.Q (result[29]), .CK (CTS_n_tid0_81), .D (n_97));
DFF_X1 \result_reg[30]  (.Q (result[30]), .CK (CTS_n_tid0_81), .D (n_98));
DFF_X1 \result_reg[31]  (.Q (result[31]), .CK (CTS_n_tid0_81), .D (n_99));
DFF_X1 \result_reg[32]  (.Q (result[32]), .CK (CTS_n_tid0_81), .D (n_100));
DFF_X1 \result_reg[33]  (.Q (result[33]), .CK (CTS_n_tid0_81), .D (n_101));
DFF_X1 \result_reg[34]  (.Q (result[34]), .CK (CTS_n_tid0_81), .D (n_102));
DFF_X1 \result_reg[35]  (.Q (result[35]), .CK (CTS_n_tid0_81), .D (n_103));
DFF_X1 \result_reg[36]  (.Q (result[36]), .CK (CTS_n_tid0_81), .D (n_104));
DFF_X1 \result_reg[37]  (.Q (result[37]), .CK (CTS_n_tid0_81), .D (n_105));
DFF_X1 \result_reg[38]  (.Q (result[38]), .CK (CTS_n_tid0_81), .D (n_106));
DFF_X1 \result_reg[39]  (.Q (result[39]), .CK (CTS_n_tid0_81), .D (n_107));
DFF_X1 \result_reg[40]  (.Q (result[40]), .CK (CTS_n_tid0_81), .D (n_108));
DFF_X1 \result_reg[41]  (.Q (result[41]), .CK (CTS_n_tid0_81), .D (n_109));
DFF_X1 \result_reg[42]  (.Q (result[42]), .CK (CTS_n_tid0_81), .D (n_110));
DFF_X1 \result_reg[43]  (.Q (result[43]), .CK (CTS_n_tid0_81), .D (n_111));
DFF_X1 \result_reg[44]  (.Q (result[44]), .CK (CTS_n_tid0_81), .D (n_112));
DFF_X1 \result_reg[45]  (.Q (result[45]), .CK (CTS_n_tid0_81), .D (n_113));
DFF_X1 \result_reg[46]  (.Q (result[46]), .CK (CTS_n_tid0_81), .D (n_114));
DFF_X1 \result_reg[47]  (.Q (result[47]), .CK (CTS_n_tid0_81), .D (n_115));
DFF_X1 \result_reg[48]  (.Q (result[48]), .CK (CTS_n_tid0_81), .D (n_116));
DFF_X1 \result_reg[49]  (.Q (result[49]), .CK (CTS_n_tid0_81), .D (n_117));
DFF_X1 \result_reg[50]  (.Q (result[50]), .CK (CTS_n_tid0_81), .D (n_118));
DFF_X1 \result_reg[51]  (.Q (result[51]), .CK (CTS_n_tid0_81), .D (n_119));
DFF_X1 \result_reg[52]  (.Q (result[52]), .CK (CTS_n_tid0_81), .D (n_120));
DFF_X1 \result_reg[53]  (.Q (result[53]), .CK (CTS_n_tid0_81), .D (n_121));
DFF_X1 \result_reg[54]  (.Q (result[54]), .CK (CTS_n_tid0_81), .D (n_122));
DFF_X1 \result_reg[55]  (.Q (result[55]), .CK (CTS_n_tid0_81), .D (n_123));
DFF_X1 \result_reg[56]  (.Q (result[56]), .CK (CTS_n_tid0_81), .D (n_124));
DFF_X1 \result_reg[57]  (.Q (result[57]), .CK (CTS_n_tid0_81), .D (n_125));
DFF_X1 \result_reg[58]  (.Q (result[58]), .CK (CTS_n_tid0_81), .D (n_126));
DFF_X1 \result_reg[59]  (.Q (result[59]), .CK (CTS_n_tid0_81), .D (n_127));
DFF_X1 \result_reg[60]  (.Q (result[60]), .CK (CTS_n_tid0_81), .D (n_128));
DFF_X1 \result_reg[61]  (.Q (result[61]), .CK (CTS_n_tid0_81), .D (n_129));
DFF_X1 \result_reg[62]  (.Q (result[62]), .CK (CTS_n_tid0_81), .D (n_130));
DFF_X1 \result_reg[63]  (.Q (result[63]), .CK (CTS_n_tid0_81), .D (n_131));
CLKGATETST_X8 clk_gate_result_reg (.GCK (CTS_n_tid0_84), .CK (CTS_n_tid0_247), .E (n_266), .SE (1'b0 ));
AOI21_X1 i_1_1137 (.ZN (n_1_938), .A (n_1_728), .B1 (n_1_704), .B2 (n_1_701));
INV_X2 i_1_1136 (.ZN (n_1_937), .A (\counter[4] ));
INV_X1 i_1_1135 (.ZN (n_1_936), .A (\counter[3] ));
INV_X2 i_1_1134 (.ZN (n_1_935), .A (\counter[2] ));
INV_X1 i_1_1133 (.ZN (n_1_934), .A (\counter[1] ));
INV_X1 i_1_1132 (.ZN (n_1_933), .A (\counter[0] ));
INV_X1 i_1_1131 (.ZN (n_1_932), .A (b[25]));
INV_X1 i_1_1130 (.ZN (n_1_931), .A (b[23]));
INV_X1 i_1_1129 (.ZN (n_1_930), .A (b[18]));
INV_X1 i_1_1128 (.ZN (n_1_929), .A (b[17]));
INV_X1 i_1_1127 (.ZN (n_1_928), .A (b[16]));
INV_X1 i_1_1126 (.ZN (n_1_927), .A (b[9]));
INV_X1 i_1_1125 (.ZN (n_1_926), .A (b[7]));
INV_X1 i_1_1124 (.ZN (n_1_925), .A (b[2]));
INV_X1 i_1_1123 (.ZN (n_1_924), .A (b[1]));
INV_X1 i_1_1122 (.ZN (n_1_923), .A (b[0]));
INV_X1 i_1_1121 (.ZN (n_1_922), .A (en));
INV_X1 i_1_1120 (.ZN (n_1_921), .A (\firstInputComplement[31] ));
INV_X1 i_1_1119 (.ZN (n_1_920), .A (\firstInputComplement[30] ));
INV_X1 i_1_1118 (.ZN (n_1_919), .A (\firstInputComplement[29] ));
INV_X1 i_1_1117 (.ZN (n_1_918), .A (\firstInputComplement[28] ));
INV_X1 i_1_1116 (.ZN (n_1_917), .A (\firstInputComplement[27] ));
INV_X1 i_1_1115 (.ZN (n_1_916), .A (\firstInputComplement[26] ));
INV_X1 i_1_1114 (.ZN (n_1_915), .A (\firstInputComplement[25] ));
INV_X1 i_1_1113 (.ZN (n_1_914), .A (\firstInputComplement[24] ));
INV_X1 i_1_1112 (.ZN (n_1_913), .A (\firstInputComplement[23] ));
INV_X1 i_1_1111 (.ZN (n_1_912), .A (\firstInputComplement[22] ));
INV_X1 i_1_1110 (.ZN (n_1_911), .A (\firstInputComplement[21] ));
INV_X1 i_1_1109 (.ZN (n_1_910), .A (\firstInputComplement[20] ));
INV_X1 i_1_1108 (.ZN (n_1_909), .A (\firstInputComplement[19] ));
INV_X1 i_1_1107 (.ZN (n_1_908), .A (\firstInputComplement[18] ));
INV_X1 i_1_1106 (.ZN (n_1_907), .A (\firstInputComplement[17] ));
INV_X1 i_1_1105 (.ZN (n_1_906), .A (\firstInputComplement[16] ));
INV_X1 i_1_1104 (.ZN (n_1_905), .A (\firstInputComplement[15] ));
INV_X1 i_1_1103 (.ZN (n_1_904), .A (\firstInputComplement[14] ));
INV_X1 i_1_1102 (.ZN (n_1_903), .A (\firstInputComplement[13] ));
INV_X1 i_1_1101 (.ZN (n_1_902), .A (\firstInputComplement[12] ));
INV_X1 i_1_1100 (.ZN (n_1_901), .A (\firstInputComplement[11] ));
INV_X1 i_1_1099 (.ZN (n_1_900), .A (\firstInputComplement[10] ));
INV_X1 i_1_1098 (.ZN (n_1_899), .A (\firstInputComplement[9] ));
INV_X1 i_1_1097 (.ZN (n_1_898), .A (\firstInputComplement[8] ));
INV_X1 i_1_1096 (.ZN (n_1_897), .A (\firstInputComplement[7] ));
INV_X1 i_1_1095 (.ZN (n_1_896), .A (\firstInputComplement[6] ));
INV_X1 i_1_1094 (.ZN (n_1_895), .A (\firstInputComplement[5] ));
INV_X1 i_1_1093 (.ZN (n_1_894), .A (\firstInputComplement[4] ));
INV_X1 i_1_1092 (.ZN (n_1_893), .A (\firstInputComplement[3] ));
INV_X1 i_1_1091 (.ZN (n_1_892), .A (\firstInputComplement[2] ));
INV_X1 i_1_1090 (.ZN (n_1_891), .A (\firstInputComplement[1] ));
INV_X1 i_1_1089 (.ZN (n_1_890), .A (a[31]));
INV_X1 i_1_1088 (.ZN (n_1_889), .A (a[30]));
INV_X1 i_1_1087 (.ZN (n_1_888), .A (a[29]));
INV_X1 i_1_1086 (.ZN (n_1_887), .A (a[28]));
INV_X1 i_1_1085 (.ZN (n_1_886), .A (a[27]));
INV_X1 i_1_1084 (.ZN (n_1_885), .A (a[26]));
INV_X1 i_1_1083 (.ZN (n_1_884), .A (a[25]));
INV_X1 i_1_1082 (.ZN (n_1_883), .A (a[24]));
INV_X1 i_1_1081 (.ZN (n_1_882), .A (a[23]));
INV_X1 i_1_1080 (.ZN (n_1_881), .A (a[22]));
INV_X1 i_1_1079 (.ZN (n_1_880), .A (a[21]));
INV_X1 i_1_1078 (.ZN (n_1_879), .A (a[20]));
INV_X1 i_1_1077 (.ZN (n_1_878), .A (a[19]));
INV_X1 i_1_1076 (.ZN (n_1_877), .A (a[18]));
INV_X1 i_1_1075 (.ZN (n_1_876), .A (a[17]));
INV_X1 i_1_1074 (.ZN (n_1_875), .A (a[16]));
INV_X1 i_1_1073 (.ZN (n_1_874), .A (a[15]));
INV_X1 i_1_1072 (.ZN (n_1_873), .A (a[14]));
INV_X1 i_1_1071 (.ZN (n_1_872), .A (a[13]));
INV_X1 i_1_1070 (.ZN (n_1_871), .A (a[12]));
INV_X1 i_1_1069 (.ZN (n_1_870), .A (a[11]));
INV_X1 i_1_1068 (.ZN (n_1_869), .A (a[10]));
INV_X1 i_1_1067 (.ZN (n_1_868), .A (a[9]));
INV_X1 i_1_1066 (.ZN (n_1_867), .A (a[8]));
INV_X1 i_1_1065 (.ZN (n_1_866), .A (a[7]));
INV_X1 i_1_1064 (.ZN (n_1_865), .A (a[6]));
INV_X1 i_1_1063 (.ZN (n_1_864), .A (a[5]));
INV_X1 i_1_1062 (.ZN (n_1_863), .A (a[4]));
INV_X1 i_1_1061 (.ZN (n_1_862), .A (a[3]));
INV_X1 i_1_1060 (.ZN (n_1_861), .A (a[2]));
INV_X1 i_1_1059 (.ZN (n_1_860), .A (a[1]));
INV_X1 i_1_1058 (.ZN (n_1_859), .A (a[0]));
INV_X1 i_1_1057 (.ZN (n_1_858), .A (n_66));
INV_X1 i_1_1056 (.ZN (n_1_857), .A (n_65));
INV_X1 i_1_1055 (.ZN (n_1_856), .A (n_64));
INV_X1 i_1_1054 (.ZN (n_1_855), .A (n_63));
INV_X1 i_1_1053 (.ZN (n_1_854), .A (n_62));
INV_X1 i_1_1052 (.ZN (n_1_853), .A (n_61));
INV_X1 i_1_1051 (.ZN (n_1_852), .A (n_60));
INV_X1 i_1_1050 (.ZN (n_1_851), .A (n_59));
INV_X1 i_1_1049 (.ZN (n_1_850), .A (n_58));
INV_X1 i_1_1048 (.ZN (n_1_849), .A (n_57));
INV_X1 i_1_1047 (.ZN (n_1_848), .A (n_56));
INV_X1 i_1_1046 (.ZN (n_1_847), .A (n_55));
INV_X1 i_1_1045 (.ZN (n_1_846), .A (n_54));
INV_X1 i_1_1044 (.ZN (n_1_845), .A (n_53));
INV_X1 i_1_1043 (.ZN (n_1_844), .A (n_52));
INV_X1 i_1_1042 (.ZN (n_1_843), .A (n_51));
INV_X1 i_1_1041 (.ZN (n_1_842), .A (n_50));
INV_X1 i_1_1040 (.ZN (n_1_841), .A (n_49));
INV_X1 i_1_1039 (.ZN (n_1_840), .A (n_48));
INV_X1 i_1_1038 (.ZN (n_1_839), .A (n_47));
INV_X1 i_1_1037 (.ZN (n_1_838), .A (n_46));
INV_X1 i_1_1036 (.ZN (n_1_837), .A (n_45));
INV_X1 i_1_1035 (.ZN (n_1_836), .A (n_44));
INV_X1 i_1_1034 (.ZN (n_1_835), .A (n_43));
INV_X1 i_1_1033 (.ZN (n_1_834), .A (n_42));
INV_X1 i_1_1032 (.ZN (n_1_833), .A (n_41));
INV_X1 i_1_1031 (.ZN (n_1_832), .A (n_40));
INV_X1 i_1_1030 (.ZN (n_1_831), .A (n_39));
INV_X1 i_1_1029 (.ZN (n_1_830), .A (n_38));
INV_X1 i_1_1028 (.ZN (n_1_829), .A (n_37));
INV_X1 i_1_1027 (.ZN (n_1_828), .A (n_36));
INV_X1 i_1_1026 (.ZN (n_1_827), .A (n_35));
INV_X1 i_1_1025 (.ZN (n_1_826), .A (n_34));
INV_X1 i_1_1024 (.ZN (n_1_825), .A (n_33));
INV_X1 i_1_1023 (.ZN (n_1_824), .A (n_32));
INV_X1 i_1_1022 (.ZN (n_1_823), .A (n_31));
INV_X1 i_1_1021 (.ZN (n_1_822), .A (n_30));
INV_X1 i_1_1020 (.ZN (n_1_821), .A (n_29));
INV_X1 i_1_1019 (.ZN (n_1_820), .A (n_28));
INV_X1 i_1_1018 (.ZN (n_1_819), .A (n_27));
INV_X1 i_1_1017 (.ZN (n_1_818), .A (n_26));
INV_X1 i_1_1016 (.ZN (n_1_817), .A (n_25));
INV_X1 i_1_1015 (.ZN (n_1_816), .A (n_24));
INV_X1 i_1_1014 (.ZN (n_1_815), .A (n_23));
INV_X1 i_1_1013 (.ZN (n_1_814), .A (n_22));
INV_X1 i_1_1012 (.ZN (n_1_813), .A (n_21));
INV_X1 i_1_1011 (.ZN (n_1_812), .A (n_20));
INV_X1 i_1_1010 (.ZN (n_1_811), .A (n_19));
INV_X1 i_1_1009 (.ZN (n_1_810), .A (n_18));
INV_X1 i_1_1008 (.ZN (n_1_809), .A (n_17));
INV_X1 i_1_1007 (.ZN (n_1_808), .A (n_16));
INV_X1 i_1_1006 (.ZN (n_1_807), .A (n_15));
INV_X1 i_1_1005 (.ZN (n_1_806), .A (n_14));
INV_X1 i_1_1004 (.ZN (n_1_805), .A (n_13));
INV_X1 i_1_1003 (.ZN (n_1_804), .A (n_12));
INV_X1 i_1_1002 (.ZN (n_1_803), .A (n_11));
INV_X1 i_1_1001 (.ZN (n_1_802), .A (n_10));
INV_X1 i_1_1000 (.ZN (n_1_801), .A (n_9));
INV_X1 i_1_999 (.ZN (n_1_800), .A (n_8));
INV_X1 i_1_998 (.ZN (n_1_799), .A (n_7));
INV_X1 i_1_997 (.ZN (n_1_798), .A (n_6));
INV_X1 i_1_996 (.ZN (n_1_797), .A (n_5));
INV_X1 i_1_995 (.ZN (n_1_796), .A (n_4));
INV_X1 i_1_994 (.ZN (n_1_795), .A (n_3));
INV_X1 i_1_993 (.ZN (n_1_794), .A (n_1_3));
INV_X1 i_1_992 (.ZN (n_1_793), .A (n_1_4));
INV_X1 i_1_991 (.ZN (n_1_792), .A (n_1_5));
XOR2_X1 i_1_990 (.Z (n_1_791), .A (n_1_937), .B (n_1_2));
NAND4_X1 i_1_989 (.ZN (n_1_790), .A1 (\counter[0] ), .A2 (n_1_794), .A3 (n_1_793), .A4 (n_1_792));
OR2_X1 i_1_988 (.ZN (n_1_789), .A1 (n_1_791), .A2 (n_1_790));
NOR2_X2 i_1_987 (.ZN (n_1_788), .A1 (\counter[1] ), .A2 (\counter[0] ));
INV_X1 i_1_986 (.ZN (n_1_787), .A (n_1_788));
NOR2_X1 i_1_985 (.ZN (n_1_786), .A1 (\counter[3] ), .A2 (\counter[2] ));
NAND3_X1 i_1_984 (.ZN (n_1_785), .A1 (n_1_788), .A2 (n_1_786), .A3 (n_1_937));
INV_X1 i_1_983 (.ZN (n_1_784), .A (hfn_ipo_n16));
OR3_X1 i_1_982 (.ZN (n_1_783), .A1 (reset), .A2 (resetReg), .A3 (hfn_ipo_n14));
OAI21_X1 i_1_981 (.ZN (n_268), .A (en), .B1 (n_1_789), .B2 (n_1_783));
OAI21_X1 i_1_980 (.ZN (n_1_782), .A (en), .B1 (reset), .B2 (resetReg));
INV_X1 i_1_979 (.ZN (n_267), .A (n_1_782));
NOR2_X1 i_1_978 (.ZN (n_1_781), .A1 (n_1_922), .A2 (hfn_ipo_n15));
OAI21_X1 i_1_977 (.ZN (n_266), .A (n_1_782), .B1 (n_1_789), .B2 (n_1_781));
NOR3_X1 i_1_976 (.ZN (n_265), .A1 (n_1_922), .A2 (reset), .A3 (resetReg));
NOR2_X1 i_1_975 (.ZN (n_1_780), .A1 (n_1_935), .A2 (n_1_933));
INV_X1 i_1_974 (.ZN (n_1_779), .A (n_1_780));
NOR2_X1 i_1_973 (.ZN (n_1_778), .A1 (n_1_936), .A2 (n_1_934));
NOR2_X2 i_1_972 (.ZN (n_1_777), .A1 (\counter[3] ), .A2 (n_1_934));
AOI22_X1 i_1_971 (.ZN (n_1_776), .A1 (b[30]), .A2 (n_1_778), .B1 (b[14]), .B2 (n_1_777));
NOR2_X1 i_1_970 (.ZN (n_1_775), .A1 (n_1_936), .A2 (\counter[1] ));
INV_X1 i_1_969 (.ZN (n_1_774), .A (n_1_775));
NOR2_X1 i_1_968 (.ZN (n_1_773), .A1 (n_1_935), .A2 (\counter[0] ));
INV_X2 i_1_967 (.ZN (n_1_772), .A (n_1_773));
AOI22_X1 i_1_966 (.ZN (n_1_771), .A1 (b[24]), .A2 (n_1_773), .B1 (b[26]), .B2 (n_1_780));
OAI22_X1 i_1_965 (.ZN (n_1_770), .A1 (n_1_779), .A2 (n_1_776), .B1 (n_1_774), .B2 (n_1_771));
AOI22_X1 i_1_964 (.ZN (n_1_769), .A1 (b[12]), .A2 (n_1_777), .B1 (b[28]), .B2 (n_1_778));
NAND2_X1 i_1_963 (.ZN (n_1_768), .A1 (n_1_936), .A2 (n_1_934));
AOI22_X1 i_1_962 (.ZN (n_1_767), .A1 (b[10]), .A2 (n_1_780), .B1 (b[8]), .B2 (n_1_773));
OAI22_X1 i_1_961 (.ZN (n_1_766), .A1 (n_1_772), .A2 (n_1_769), .B1 (n_1_768), .B2 (n_1_767));
NOR2_X1 i_1_960 (.ZN (n_1_765), .A1 (n_1_770), .A2 (n_1_766));
NOR2_X1 i_1_959 (.ZN (n_1_764), .A1 (\counter[2] ), .A2 (n_1_933));
INV_X1 i_1_958 (.ZN (n_1_763), .A (n_1_764));
OAI22_X1 i_1_957 (.ZN (n_1_762), .A1 (n_1_930), .A2 (n_1_774), .B1 (n_1_925), .B2 (n_1_768));
AOI221_X1 i_1_956 (.ZN (n_1_761), .A (n_1_762), .B1 (b[6]), .B2 (n_1_777), .C1 (b[22]), .C2 (n_1_778));
NAND2_X1 i_1_955 (.ZN (n_1_760), .A1 (n_1_935), .A2 (n_1_933));
OAI22_X1 i_1_954 (.ZN (n_1_759), .A1 (n_1_923), .A2 (n_1_768), .B1 (n_1_928), .B2 (n_1_774));
AOI221_X1 i_1_953 (.ZN (n_1_758), .A (n_1_759), .B1 (b[20]), .B2 (n_1_778), .C1 (b[4]), .C2 (n_1_777));
OAI221_X1 i_1_952 (.ZN (n_1_757), .A (n_1_765), .B1 (n_1_763), .B2 (n_1_761), .C1 (n_1_760), .C2 (n_1_758));
AOI222_X1 i_1_951 (.ZN (n_1_756), .A1 (b[3]), .A2 (n_1_777), .B1 (b[15]), .B2 (n_1_775)
    , .C1 (b[19]), .C2 (n_1_778));
OAI22_X1 i_1_950 (.ZN (n_1_755), .A1 (n_1_927), .A2 (n_1_768), .B1 (n_1_932), .B2 (n_1_774));
AOI221_X1 i_1_949 (.ZN (n_1_754), .A (n_1_755), .B1 (b[29]), .B2 (n_1_778), .C1 (b[13]), .C2 (n_1_777));
OAI22_X1 i_1_948 (.ZN (n_1_753), .A1 (n_1_760), .A2 (n_1_756), .B1 (n_1_779), .B2 (n_1_754));
INV_X1 i_1_947 (.ZN (n_1_752), .A (n_1_753));
OAI22_X1 i_1_946 (.ZN (n_1_751), .A1 (n_1_924), .A2 (n_1_768), .B1 (n_1_929), .B2 (n_1_774));
AOI221_X1 i_1_945 (.ZN (n_1_750), .A (n_1_751), .B1 (b[5]), .B2 (n_1_777), .C1 (b[21]), .C2 (n_1_778));
OAI22_X1 i_1_944 (.ZN (n_1_749), .A1 (n_1_931), .A2 (n_1_774), .B1 (n_1_926), .B2 (n_1_768));
AOI221_X1 i_1_943 (.ZN (n_1_748), .A (n_1_749), .B1 (b[11]), .B2 (n_1_777), .C1 (b[27]), .C2 (n_1_778));
OAI221_X1 i_1_942 (.ZN (n_1_747), .A (n_1_752), .B1 (n_1_763), .B2 (n_1_750), .C1 (n_1_772), .C2 (n_1_748));
NAND2_X1 i_1_941 (.ZN (n_1_746), .A1 (n_1_757), .A2 (n_1_747));
OR2_X1 i_1_940 (.ZN (n_1_745), .A1 (n_1_757), .A2 (n_1_747));
NAND2_X1 i_1_939 (.ZN (n_1_744), .A1 (n_1_746), .A2 (n_1_745));
AOI22_X1 i_1_938 (.ZN (n_1_743), .A1 (b[23]), .A2 (n_1_778), .B1 (b[7]), .B2 (n_1_777));
AOI22_X1 i_1_937 (.ZN (n_1_742), .A1 (b[15]), .A2 (n_1_777), .B1 (b[31]), .B2 (n_1_778));
OAI22_X1 i_1_936 (.ZN (n_1_741), .A1 (n_1_763), .A2 (n_1_743), .B1 (n_1_779), .B2 (n_1_742));
AOI22_X1 i_1_935 (.ZN (n_1_740), .A1 (b[19]), .A2 (n_1_764), .B1 (b[27]), .B2 (n_1_780));
AOI22_X1 i_1_934 (.ZN (n_1_739), .A1 (b[11]), .A2 (n_1_780), .B1 (b[3]), .B2 (n_1_764));
OAI22_X1 i_1_933 (.ZN (n_1_738), .A1 (n_1_774), .A2 (n_1_740), .B1 (n_1_768), .B2 (n_1_739));
OAI22_X1 i_1_932 (.ZN (n_1_737), .A1 (n_1_760), .A2 (n_1_750), .B1 (n_1_772), .B2 (n_1_754));
NOR3_X1 i_1_931 (.ZN (n_1_736), .A1 (n_1_741), .A2 (n_1_738), .A3 (n_1_737));
INV_X1 i_1_930 (.ZN (n_1_735), .A (n_1_736));
OR2_X2 i_1_929 (.ZN (n_1_734), .A1 (n_1_744), .A2 (n_1_736));
OR2_X2 i_1_928 (.ZN (n_1_733), .A1 (n_1_744), .A2 (n_1_735));
NOR2_X4 i_1_927 (.ZN (n_1_732), .A1 (n_1_746), .A2 (n_1_735));
NOR2_X4 i_1_926 (.ZN (n_1_731), .A1 (n_1_745), .A2 (n_1_736));
AOI22_X1 i_1_925 (.ZN (n_1_730), .A1 (a[30]), .A2 (n_1_732), .B1 (\firstInputComplement[30] ), .B2 (n_1_731));
OAI221_X1 i_1_924 (.ZN (n_1_729), .A (n_1_730), .B1 (n_1_890), .B2 (n_1_733), .C1 (n_1_921), .C2 (n_1_734));
INV_X1 i_1_923 (.ZN (n_1_728), .A (n_1_729));
NAND3_X1 i_1_922 (.ZN (n_1_727), .A1 (n_1_935), .A2 (n_1_933), .A3 (\counter[1] ));
NAND2_X1 i_1_921 (.ZN (n_1_726), .A1 (n_1_937), .A2 (\counter[3] ));
NOR2_X1 i_1_920 (.ZN (n_1_725), .A1 (n_1_727), .A2 (n_1_726));
INV_X2 i_1_919 (.ZN (n_1_724), .A (n_1_725));
NOR2_X1 i_1_918 (.ZN (n_1_723), .A1 (n_1_728), .A2 (n_1_724));
NAND2_X1 i_1_917 (.ZN (n_1_722), .A1 (n_1_937), .A2 (n_1_936));
NAND3_X1 i_1_916 (.ZN (n_1_721), .A1 (n_1_937), .A2 (n_1_936), .A3 (n_1_729));
OR2_X1 i_1_915 (.ZN (n_1_720), .A1 (n_1_934), .A2 (n_1_721));
NOR2_X1 i_1_914 (.ZN (n_1_719), .A1 (n_1_773), .A2 (n_1_720));
OR2_X1 i_1_913 (.ZN (n_1_718), .A1 (n_1_723), .A2 (n_1_719));
NAND2_X1 i_1_912 (.ZN (n_1_717), .A1 (\counter[1] ), .A2 (\counter[0] ));
NAND3_X1 i_1_911 (.ZN (n_1_716), .A1 (\counter[1] ), .A2 (\counter[0] ), .A3 (\counter[2] ));
NOR2_X1 i_1_910 (.ZN (n_1_715), .A1 (n_1_935), .A2 (n_1_934));
INV_X1 i_1_909 (.ZN (n_1_714), .A (n_1_715));
NAND4_X2 i_1_908 (.ZN (n_1_713), .A1 (n_1_936), .A2 (n_1_716), .A3 (n_1_937), .A4 (n_1_715));
INV_X1 i_1_907 (.ZN (n_1_712), .A (n_1_713));
NOR2_X1 i_1_906 (.ZN (n_1_711), .A1 (n_1_728), .A2 (n_1_713));
INV_X1 i_1_905 (.ZN (n_1_710), .A (n_1_711));
NAND3_X1 i_1_904 (.ZN (n_1_709), .A1 (n_1_937), .A2 (n_1_936), .A3 (n_1_934));
NOR2_X2 i_1_903 (.ZN (n_1_708), .A1 (n_1_779), .A2 (n_1_709));
INV_X1 i_1_902 (.ZN (n_1_707), .A (n_1_708));
NOR2_X1 i_1_901 (.ZN (n_1_706), .A1 (n_1_728), .A2 (n_1_707));
OAI21_X1 i_1_900 (.ZN (n_1_705), .A (n_1_710), .B1 (n_1_728), .B2 (n_1_707));
NAND4_X4 i_1_899 (.ZN (n_1_704), .A1 (n_1_937), .A2 (\counter[3] ), .A3 (n_1_935), .A4 (n_1_788));
NOR2_X1 i_1_898 (.ZN (n_1_703), .A1 (n_1_728), .A2 (n_1_704));
NOR3_X1 i_1_897 (.ZN (n_1_702), .A1 (n_1_774), .A2 (n_1_763), .A3 (\counter[4] ));
INV_X2 i_1_896 (.ZN (n_1_701), .A (n_1_702));
OR2_X1 i_1_895 (.ZN (n_1_700), .A1 (n_1_705), .A2 (n_1_938));
NOR2_X1 i_1_894 (.ZN (n_1_699), .A1 (hfn_ipo_n15), .A2 (n_1_728));
INV_X1 i_1_893 (.ZN (n_1_698), .A (n_1_699));
NOR2_X1 i_1_892 (.ZN (n_1_697), .A1 (n_1_763), .A2 (n_1_709));
INV_X1 i_1_891 (.ZN (n_1_696), .A (n_1_697));
NOR2_X1 i_1_890 (.ZN (n_1_695), .A1 (n_1_728), .A2 (n_1_696));
NOR2_X1 i_1_889 (.ZN (n_1_694), .A1 (n_1_699), .A2 (n_1_695));
INV_X1 i_1_888 (.ZN (n_1_693), .A (n_1_694));
OR2_X4 i_1_887 (.ZN (n_1_692), .A1 (n_1_772), .A2 (n_1_709));
NOR2_X1 i_1_886 (.ZN (n_1_691), .A1 (n_1_728), .A2 (n_1_692));
OAI21_X1 i_1_885 (.ZN (n_1_690), .A (n_1_694), .B1 (n_1_728), .B2 (n_1_692));
NOR2_X1 i_1_884 (.ZN (n_1_689), .A1 (n_1_700), .A2 (n_1_690));
OR3_X1 i_1_883 (.ZN (n_1_688), .A1 (n_1_700), .A2 (n_1_690), .A3 (n_1_718));
OR4_X1 i_1_882 (.ZN (n_1_687), .A1 (n_1_774), .A2 (n_1_763), .A3 (n_1_937), .A4 (n_1_786));
AOI22_X1 i_1_881 (.ZN (n_1_686), .A1 (a[12]), .A2 (n_1_732), .B1 (\firstInputComplement[12] ), .B2 (n_1_731));
OAI221_X1 i_1_880 (.ZN (n_1_685), .A (n_1_686), .B1 (n_1_872), .B2 (n_1_733), .C1 (n_1_903), .C2 (n_1_734));
INV_X1 i_1_879 (.ZN (n_1_684), .A (n_1_685));
NAND2_X1 i_1_878 (.ZN (n_1_683), .A1 (\counter[4] ), .A2 (\counter[3] ));
NOR2_X1 i_1_877 (.ZN (n_1_682), .A1 (n_1_714), .A2 (n_1_683));
NAND2_X1 i_1_876 (.ZN (n_1_681), .A1 (n_1_717), .A2 (n_1_682));
AOI22_X1 i_1_875 (.ZN (n_1_680), .A1 (a[2]), .A2 (n_1_732), .B1 (\firstInputComplement[2] ), .B2 (n_1_731));
OAI221_X2 i_1_874 (.ZN (n_1_679), .A (n_1_680), .B1 (n_1_862), .B2 (n_1_733), .C1 (n_1_893), .C2 (n_1_734));
INV_X2 i_1_873 (.ZN (n_1_678), .A (n_1_679));
NAND2_X1 i_1_872 (.ZN (n_1_677), .A1 (\counter[0] ), .A2 (n_1_682));
OAI21_X1 i_1_871 (.ZN (n_1_676), .A (a[0]), .B1 (n_1_732), .B2 (n_1_731));
OAI221_X1 i_1_870 (.ZN (n_1_675), .A (n_1_676), .B1 (n_1_891), .B2 (n_1_734), .C1 (n_1_860), .C2 (n_1_733));
INV_X2 i_1_869 (.ZN (n_1_674), .A (n_1_675));
NAND3_X2 i_1_868 (.ZN (n_1_673), .A1 (\counter[4] ), .A2 (n_1_780), .A3 (n_1_777));
AOI22_X1 i_1_867 (.ZN (n_1_672), .A1 (a[16]), .A2 (n_1_732), .B1 (\firstInputComplement[16] ), .B2 (n_1_731));
OAI221_X1 i_1_866 (.ZN (n_1_671), .A (n_1_672), .B1 (n_1_876), .B2 (n_1_733), .C1 (n_1_907), .C2 (n_1_734));
INV_X2 i_1_865 (.ZN (n_1_670), .A (n_1_671));
OAI22_X1 i_1_864 (.ZN (n_1_669), .A1 (n_1_677), .A2 (n_1_674), .B1 (n_1_673), .B2 (n_1_670));
NOR3_X1 i_1_863 (.ZN (n_1_668), .A1 (n_1_935), .A2 (n_1_787), .A3 (n_1_683));
INV_X1 i_1_862 (.ZN (n_1_667), .A (n_1_668));
AOI22_X1 i_1_861 (.ZN (n_1_666), .A1 (a[6]), .A2 (n_1_732), .B1 (\firstInputComplement[6] ), .B2 (n_1_731));
OAI221_X1 i_1_860 (.ZN (n_1_665), .A (n_1_666), .B1 (n_1_866), .B2 (n_1_733), .C1 (n_1_897), .C2 (n_1_734));
INV_X1 i_1_859 (.ZN (n_1_664), .A (drc_ipo_n19));
NAND2_X1 i_1_858 (.ZN (n_1_663), .A1 (n_1_937), .A2 (n_1_778));
NOR2_X2 i_1_857 (.ZN (n_1_662), .A1 (n_1_763), .A2 (n_1_663));
INV_X1 i_1_856 (.ZN (n_1_661), .A (n_1_662));
NOR2_X1 i_1_855 (.ZN (n_1_660), .A1 (n_1_728), .A2 (n_1_661));
AOI211_X1 i_1_854 (.ZN (n_1_659), .A (n_1_660), .B (n_1_669), .C1 (n_1_668), .C2 (drc_ipo_n19));
OAI221_X1 i_1_853 (.ZN (n_1_658), .A (n_1_659), .B1 (n_1_687), .B2 (n_1_684), .C1 (n_1_681), .C2 (n_1_678));
NOR4_X1 i_1_852 (.ZN (n_1_657), .A1 (\counter[3] ), .A2 (\counter[2] ), .A3 (n_1_937), .A4 (\counter[1] ));
NAND2_X2 i_1_851 (.ZN (n_1_656), .A1 (\counter[0] ), .A2 (n_1_657));
AOI22_X1 i_1_850 (.ZN (n_1_655), .A1 (a[28]), .A2 (n_1_732), .B1 (\firstInputComplement[28] ), .B2 (n_1_731));
OAI221_X1 i_1_849 (.ZN (n_1_654), .A (n_1_655), .B1 (n_1_888), .B2 (n_1_733), .C1 (n_1_919), .C2 (n_1_734));
INV_X1 i_1_848 (.ZN (n_1_653), .A (n_1_654));
OR3_X1 i_1_847 (.ZN (n_1_652), .A1 (\counter[2] ), .A2 (n_1_717), .A3 (n_1_683));
AOI22_X1 i_1_846 (.ZN (n_1_651), .A1 (a[8]), .A2 (n_1_732), .B1 (\firstInputComplement[8] ), .B2 (n_1_731));
OAI221_X1 i_1_845 (.ZN (n_1_650), .A (n_1_651), .B1 (n_1_868), .B2 (n_1_733), .C1 (n_1_899), .C2 (n_1_734));
INV_X2 i_1_844 (.ZN (n_1_649), .A (n_1_650));
NOR3_X4 i_1_843 (.ZN (n_1_648), .A1 (\counter[4] ), .A2 (n_1_774), .A3 (n_1_779));
INV_X1 i_1_842 (.ZN (n_1_647), .A (n_1_648));
NOR3_X2 i_1_841 (.ZN (n_1_646), .A1 (n_1_935), .A2 (n_1_787), .A3 (n_1_726));
INV_X2 i_1_840 (.ZN (n_1_645), .A (n_1_646));
NAND2_X1 i_1_839 (.ZN (n_1_644), .A1 (n_1_647), .A2 (n_1_645));
NOR3_X1 i_1_838 (.ZN (n_1_643), .A1 (\counter[4] ), .A2 (n_1_714), .A3 (n_1_936));
OAI21_X1 i_1_837 (.ZN (n_1_642), .A (n_1_729), .B1 (n_1_644), .B2 (n_1_643));
NAND3_X1 i_1_836 (.ZN (n_1_641), .A1 (\counter[4] ), .A2 (n_1_786), .A3 (\counter[1] ));
OR2_X1 i_1_835 (.ZN (n_1_640), .A1 (n_1_933), .A2 (n_1_641));
AOI22_X1 i_1_834 (.ZN (n_1_639), .A1 (a[24]), .A2 (n_1_732), .B1 (\firstInputComplement[24] ), .B2 (n_1_731));
OAI221_X1 i_1_833 (.ZN (n_1_638), .A (n_1_639), .B1 (n_1_884), .B2 (n_1_733), .C1 (n_1_915), .C2 (n_1_734));
INV_X1 i_1_832 (.ZN (n_1_637), .A (n_1_638));
OAI21_X1 i_1_831 (.ZN (n_1_636), .A (n_1_642), .B1 (CLOCK_sgo__n273), .B2 (n_1_637));
INV_X1 i_1_830 (.ZN (n_1_635), .A (n_1_636));
OAI221_X1 i_1_829 (.ZN (n_1_634), .A (n_1_635), .B1 (n_1_656), .B2 (n_1_653), .C1 (n_1_652), .C2 (n_1_649));
NOR3_X2 i_1_828 (.ZN (n_1_633), .A1 (\counter[2] ), .A2 (n_1_787), .A3 (n_1_683));
INV_X1 i_1_827 (.ZN (n_1_632), .A (n_1_633));
AOI22_X1 i_1_826 (.ZN (n_1_631), .A1 (a[14]), .A2 (n_1_732), .B1 (\firstInputComplement[14] ), .B2 (n_1_731));
OAI221_X1 i_1_825 (.ZN (n_1_630), .A (n_1_631), .B1 (n_1_874), .B2 (n_1_733), .C1 (n_1_905), .C2 (n_1_734));
INV_X2 i_1_824 (.ZN (n_1_629), .A (n_1_630));
OR2_X1 i_1_823 (.ZN (n_1_628), .A1 (n_1_727), .A2 (n_1_683));
AOI22_X1 i_1_822 (.ZN (n_1_627), .A1 (a[10]), .A2 (n_1_732), .B1 (\firstInputComplement[10] ), .B2 (n_1_731));
OAI221_X1 i_1_821 (.ZN (n_1_626), .A (n_1_627), .B1 (n_1_870), .B2 (n_1_733), .C1 (n_1_901), .C2 (n_1_734));
INV_X2 i_1_820 (.ZN (n_1_625), .A (n_1_626));
OAI22_X1 i_1_819 (.ZN (n_1_624), .A1 (n_1_632), .A2 (n_1_629), .B1 (n_1_628), .B2 (n_1_625));
INV_X1 i_1_818 (.ZN (n_1_623), .A (n_1_624));
NOR2_X1 i_1_817 (.ZN (n_1_622), .A1 (\counter[0] ), .A2 (n_1_641));
INV_X2 i_1_816 (.ZN (n_1_621), .A (n_1_622));
AOI22_X1 i_1_815 (.ZN (n_1_620), .A1 (a[26]), .A2 (n_1_732), .B1 (\firstInputComplement[26] ), .B2 (n_1_731));
OAI221_X1 i_1_814 (.ZN (n_1_619), .A (n_1_620), .B1 (n_1_886), .B2 (n_1_733), .C1 (n_1_917), .C2 (n_1_734));
INV_X1 i_1_813 (.ZN (n_1_618), .A (n_1_619));
NAND3_X2 i_1_812 (.ZN (n_1_617), .A1 (\counter[4] ), .A2 (n_1_786), .A3 (n_1_788));
INV_X1 i_1_811 (.ZN (n_1_616), .A (n_1_617));
OAI221_X1 i_1_810 (.ZN (n_1_615), .A (n_1_623), .B1 (n_1_621), .B2 (n_1_618), .C1 (n_1_728), .C2 (n_1_617));
OAI21_X1 i_1_809 (.ZN (n_1_614), .A (n_1_936), .B1 (n_1_935), .B2 (n_1_788));
NAND4_X1 i_1_808 (.ZN (n_1_613), .A1 (n_1_936), .A2 (n_1_716), .A3 (\counter[4] ), .A4 (n_1_614));
OR2_X2 i_1_807 (.ZN (n_1_612), .A1 (n_1_715), .A2 (n_1_613));
AOI22_X1 i_1_806 (.ZN (n_1_611), .A1 (a[20]), .A2 (n_1_732), .B1 (\firstInputComplement[20] ), .B2 (n_1_731));
OAI221_X1 i_1_805 (.ZN (n_1_610), .A (n_1_611), .B1 (n_1_880), .B2 (n_1_733), .C1 (n_1_911), .C2 (n_1_734));
INV_X1 i_1_804 (.ZN (n_1_609), .A (n_1_610));
OR3_X2 i_1_803 (.ZN (n_1_608), .A1 (n_1_937), .A2 (n_1_786), .A3 (n_1_614));
AOI22_X1 i_1_802 (.ZN (n_1_607), .A1 (a[22]), .A2 (n_1_732), .B1 (\firstInputComplement[22] ), .B2 (n_1_731));
OAI221_X1 i_1_801 (.ZN (n_1_606), .A (n_1_607), .B1 (n_1_882), .B2 (n_1_733), .C1 (n_1_913), .C2 (n_1_734));
INV_X1 i_1_800 (.ZN (n_1_605), .A (n_1_606));
OAI22_X1 i_1_799 (.ZN (n_1_604), .A1 (n_1_612), .A2 (n_1_609), .B1 (n_1_608), .B2 (n_1_605));
OR4_X1 i_1_798 (.ZN (n_1_603), .A1 (n_1_935), .A2 (n_1_788), .A3 (n_1_715), .A4 (n_1_683));
AOI22_X1 i_1_797 (.ZN (n_1_602), .A1 (a[4]), .A2 (n_1_732), .B1 (\firstInputComplement[4] ), .B2 (n_1_731));
OAI221_X2 i_1_796 (.ZN (n_1_601), .A (n_1_602), .B1 (n_1_864), .B2 (n_1_733), .C1 (n_1_895), .C2 (n_1_734));
INV_X2 i_1_795 (.ZN (n_1_600), .A (n_1_601));
OR2_X1 i_1_794 (.ZN (n_1_599), .A1 (n_1_714), .A2 (n_1_613));
AOI22_X1 i_1_793 (.ZN (n_1_598), .A1 (a[18]), .A2 (n_1_732), .B1 (\firstInputComplement[18] ), .B2 (n_1_731));
OAI221_X1 i_1_792 (.ZN (n_1_597), .A (n_1_598), .B1 (n_1_878), .B2 (n_1_733), .C1 (n_1_909), .C2 (n_1_734));
INV_X1 i_1_791 (.ZN (n_1_596), .A (n_1_597));
OAI22_X1 i_1_790 (.ZN (n_1_595), .A1 (n_1_603), .A2 (n_1_600), .B1 (n_1_599), .B2 (n_1_596));
OR4_X1 i_1_789 (.ZN (n_1_594), .A1 (n_1_604), .A2 (n_1_595), .A3 (n_1_615), .A4 (n_1_634));
OR3_X1 i_1_788 (.ZN (n_264), .A1 (n_1_658), .A2 (n_1_594), .A3 (n_1_688));
NOR2_X1 i_1_787 (.ZN (n_1_593), .A1 (\counter[2] ), .A2 (n_1_720));
OAI21_X1 i_1_786 (.ZN (n_1_592), .A (n_1_694), .B1 (\counter[2] ), .B2 (n_1_720));
OR2_X1 i_1_785 (.ZN (n_1_591), .A1 (n_1_691), .A2 (n_1_592));
NOR2_X1 i_1_784 (.ZN (n_1_590), .A1 (n_1_721), .A2 (n_1_716));
OR2_X1 i_1_783 (.ZN (n_1_589), .A1 (n_1_705), .A2 (n_1_590));
OR2_X1 i_1_782 (.ZN (n_1_588), .A1 (n_1_591), .A2 (n_1_589));
OR2_X1 i_1_781 (.ZN (n_1_587), .A1 (n_1_723), .A2 (n_1_660));
OR2_X1 i_1_780 (.ZN (n_1_586), .A1 (n_1_938), .A2 (n_1_587));
OR2_X1 i_1_779 (.ZN (n_1_585), .A1 (n_1_588), .A2 (n_1_586));
OR2_X2 i_1_778 (.ZN (n_1_584), .A1 (n_1_859), .A2 (n_1_744));
AOI22_X1 i_1_777 (.ZN (n_1_583), .A1 (a[13]), .A2 (n_1_732), .B1 (\firstInputComplement[13] ), .B2 (n_1_731));
OAI221_X2 i_1_776 (.ZN (n_1_582), .A (n_1_583), .B1 (n_1_873), .B2 (n_1_733), .C1 (n_1_904), .C2 (n_1_734));
INV_X1 i_1_775 (.ZN (n_1_581), .A (n_1_582));
AOI22_X1 i_1_774 (.ZN (n_1_580), .A1 (a[5]), .A2 (n_1_732), .B1 (\firstInputComplement[5] ), .B2 (n_1_731));
OAI221_X2 i_1_773 (.ZN (n_1_579), .A (n_1_580), .B1 (n_1_865), .B2 (n_1_733), .C1 (n_1_896), .C2 (n_1_734));
INV_X2 i_1_772 (.ZN (n_1_578), .A (n_1_579));
AOI22_X1 i_1_771 (.ZN (n_1_577), .A1 (a[3]), .A2 (n_1_732), .B1 (\firstInputComplement[3] ), .B2 (n_1_731));
OAI221_X2 i_1_770 (.ZN (n_1_576), .A (n_1_577), .B1 (n_1_863), .B2 (n_1_733), .C1 (n_1_894), .C2 (n_1_734));
INV_X1 i_1_769 (.ZN (n_1_575), .A (n_1_576));
AOI22_X1 i_1_768 (.ZN (n_1_574), .A1 (a[27]), .A2 (n_1_732), .B1 (\firstInputComplement[27] ), .B2 (n_1_731));
OAI221_X1 i_1_767 (.ZN (n_1_573), .A (n_1_574), .B1 (n_1_887), .B2 (n_1_733), .C1 (n_1_918), .C2 (n_1_734));
INV_X1 i_1_766 (.ZN (n_1_572), .A (n_1_573));
OAI22_X1 i_1_765 (.ZN (n_1_571), .A1 (n_1_603), .A2 (n_1_575), .B1 (n_1_656), .B2 (n_1_572));
AOI221_X1 i_1_764 (.ZN (n_1_570), .A (n_1_571), .B1 (n_1_633), .B2 (n_1_582), .C1 (n_1_668), .C2 (n_1_579));
OAI211_X1 i_1_763 (.ZN (n_1_569), .A (n_1_642), .B (n_1_570), .C1 (n_1_677), .C2 (n_1_584));
AOI22_X1 i_1_762 (.ZN (n_1_568), .A1 (a[17]), .A2 (n_1_732), .B1 (\firstInputComplement[17] ), .B2 (n_1_731));
OAI221_X1 i_1_761 (.ZN (n_1_567), .A (n_1_568), .B1 (n_1_877), .B2 (n_1_733), .C1 (n_1_908), .C2 (n_1_734));
INV_X1 i_1_760 (.ZN (n_1_566), .A (n_1_567));
AOI22_X1 i_1_759 (.ZN (n_1_565), .A1 (a[29]), .A2 (n_1_732), .B1 (\firstInputComplement[29] ), .B2 (n_1_731));
OAI221_X1 i_1_758 (.ZN (n_1_564), .A (n_1_565), .B1 (n_1_889), .B2 (n_1_733), .C1 (n_1_920), .C2 (n_1_734));
INV_X1 i_1_757 (.ZN (n_1_563), .A (n_1_564));
AOI22_X1 i_1_756 (.ZN (n_1_562), .A1 (a[25]), .A2 (n_1_732), .B1 (\firstInputComplement[25] ), .B2 (n_1_731));
OAI221_X1 i_1_755 (.ZN (n_1_561), .A (n_1_562), .B1 (n_1_885), .B2 (n_1_733), .C1 (n_1_916), .C2 (n_1_734));
INV_X1 i_1_754 (.ZN (n_1_560), .A (n_1_561));
OAI222_X1 i_1_753 (.ZN (n_1_559), .A1 (n_1_617), .A2 (n_1_563), .B1 (n_1_621), .B2 (n_1_560)
    , .C1 (n_1_599), .C2 (n_1_566));
AOI22_X1 i_1_752 (.ZN (n_1_558), .A1 (a[23]), .A2 (n_1_732), .B1 (\firstInputComplement[23] ), .B2 (n_1_731));
OAI221_X1 i_1_751 (.ZN (n_1_557), .A (n_1_558), .B1 (n_1_883), .B2 (n_1_733), .C1 (n_1_914), .C2 (n_1_734));
INV_X1 i_1_750 (.ZN (n_1_556), .A (n_1_557));
AOI22_X1 i_1_749 (.ZN (n_1_555), .A1 (a[21]), .A2 (n_1_732), .B1 (\firstInputComplement[21] ), .B2 (n_1_731));
OAI221_X1 i_1_748 (.ZN (n_1_554), .A (n_1_555), .B1 (n_1_881), .B2 (n_1_733), .C1 (n_1_912), .C2 (n_1_734));
INV_X1 i_1_747 (.ZN (n_1_553), .A (n_1_554));
AOI22_X1 i_1_746 (.ZN (n_1_552), .A1 (a[15]), .A2 (n_1_732), .B1 (\firstInputComplement[15] ), .B2 (n_1_731));
OAI221_X1 i_1_745 (.ZN (n_1_551), .A (n_1_552), .B1 (n_1_875), .B2 (n_1_733), .C1 (n_1_906), .C2 (n_1_734));
INV_X1 i_1_744 (.ZN (n_1_550), .A (n_1_551));
AOI22_X1 i_1_743 (.ZN (n_1_549), .A1 (a[9]), .A2 (n_1_732), .B1 (\firstInputComplement[9] ), .B2 (n_1_731));
OAI221_X2 i_1_742 (.ZN (n_1_548), .A (n_1_549), .B1 (n_1_869), .B2 (n_1_733), .C1 (n_1_900), .C2 (n_1_734));
INV_X2 i_1_741 (.ZN (n_1_547), .A (n_1_548));
OAI22_X1 i_1_740 (.ZN (n_1_546), .A1 (n_1_673), .A2 (n_1_550), .B1 (n_1_628), .B2 (n_1_547));
INV_X1 i_1_739 (.ZN (n_1_545), .A (n_1_546));
OAI221_X1 i_1_738 (.ZN (n_1_544), .A (n_1_545), .B1 (CLOCK_sgo__n273), .B2 (n_1_556)
    , .C1 (n_1_608), .C2 (n_1_553));
AOI22_X1 i_1_737 (.ZN (n_1_543), .A1 (a[11]), .A2 (n_1_732), .B1 (\firstInputComplement[11] ), .B2 (n_1_731));
OAI221_X2 i_1_736 (.ZN (n_1_542), .A (n_1_543), .B1 (n_1_871), .B2 (n_1_733), .C1 (n_1_902), .C2 (n_1_734));
INV_X1 i_1_735 (.ZN (n_1_541), .A (n_1_542));
AOI22_X1 i_1_734 (.ZN (n_1_540), .A1 (a[19]), .A2 (n_1_732), .B1 (\firstInputComplement[19] ), .B2 (n_1_731));
OAI221_X1 i_1_733 (.ZN (n_1_539), .A (n_1_540), .B1 (n_1_879), .B2 (n_1_733), .C1 (n_1_910), .C2 (n_1_734));
INV_X1 i_1_732 (.ZN (n_1_538), .A (n_1_539));
OAI22_X1 i_1_731 (.ZN (n_1_537), .A1 (n_1_687), .A2 (n_1_541), .B1 (n_1_612), .B2 (n_1_538));
AOI22_X1 i_1_730 (.ZN (n_1_536), .A1 (a[7]), .A2 (n_1_732), .B1 (\firstInputComplement[7] ), .B2 (n_1_731));
OAI221_X2 i_1_729 (.ZN (n_1_535), .A (n_1_536), .B1 (n_1_867), .B2 (n_1_733), .C1 (n_1_898), .C2 (n_1_734));
INV_X1 i_1_728 (.ZN (n_1_534), .A (n_1_535));
AOI22_X1 i_1_727 (.ZN (n_1_533), .A1 (a[1]), .A2 (n_1_732), .B1 (\firstInputComplement[1] ), .B2 (n_1_731));
OAI221_X2 i_1_726 (.ZN (n_1_532), .A (n_1_533), .B1 (n_1_861), .B2 (n_1_733), .C1 (n_1_892), .C2 (n_1_734));
INV_X2 i_1_725 (.ZN (n_1_531), .A (n_1_532));
OAI22_X1 i_1_724 (.ZN (n_1_530), .A1 (n_1_652), .A2 (n_1_534), .B1 (n_1_681), .B2 (n_1_531));
OR4_X1 i_1_723 (.ZN (n_1_529), .A1 (n_1_537), .A2 (n_1_530), .A3 (n_1_544), .A4 (n_1_559));
OR3_X1 i_1_722 (.ZN (n_263), .A1 (n_1_569), .A2 (n_1_529), .A3 (n_1_585));
OAI22_X1 i_1_721 (.ZN (n_1_528), .A1 (n_1_653), .A2 (n_1_617), .B1 (n_1_637), .B2 (n_1_621));
OAI22_X1 i_1_720 (.ZN (n_1_527), .A1 (n_1_649), .A2 (n_1_628), .B1 (n_1_612), .B2 (n_1_596));
OAI21_X1 i_1_719 (.ZN (n_1_526), .A (n_1_642), .B1 (n_1_609), .B2 (n_1_608));
OAI22_X1 i_1_718 (.ZN (n_1_525), .A1 (n_1_667), .A2 (n_1_600), .B1 (n_1_670), .B2 (n_1_599));
OR4_X1 i_1_717 (.ZN (n_1_524), .A1 (n_1_528), .A2 (n_1_527), .A3 (n_1_526), .A4 (n_1_525));
OAI22_X1 i_1_716 (.ZN (n_1_523), .A1 (n_1_673), .A2 (n_1_629), .B1 (CLOCK_sgo__n273), .B2 (n_1_605));
INV_X1 i_1_715 (.ZN (n_1_522), .A (n_1_523));
OAI221_X1 i_1_714 (.ZN (n_1_521), .A (n_1_522), .B1 (n_1_684), .B2 (n_1_632), .C1 (n_1_656), .C2 (n_1_618));
OAI22_X1 i_1_713 (.ZN (n_1_520), .A1 (n_1_681), .A2 (n_1_674), .B1 (n_1_664), .B2 (n_1_652));
INV_X1 i_1_712 (.ZN (n_1_519), .A (n_1_520));
OAI221_X1 i_1_711 (.ZN (n_1_518), .A (n_1_519), .B1 (n_1_678), .B2 (n_1_603), .C1 (n_1_687), .C2 (n_1_625));
OR4_X1 i_1_710 (.ZN (n_262), .A1 (n_1_521), .A2 (n_1_518), .A3 (n_1_524), .A4 (n_1_585));
NOR2_X1 i_1_709 (.ZN (n_1_517), .A1 (n_1_772), .A2 (n_1_663));
INV_X2 i_1_708 (.ZN (n_1_516), .A (n_1_517));
NOR3_X1 i_1_707 (.ZN (n_1_515), .A1 (n_1_662), .A2 (n_1_517), .A3 (n_1_644));
OAI21_X1 i_1_706 (.ZN (n_1_514), .A (n_1_689), .B1 (n_1_728), .B2 (n_1_515));
OAI22_X1 i_1_705 (.ZN (n_1_513), .A1 (n_1_667), .A2 (n_1_575), .B1 (n_1_628), .B2 (n_1_534));
INV_X1 i_1_704 (.ZN (n_1_512), .A (n_1_513));
OAI221_X1 i_1_703 (.ZN (n_1_511), .A (n_1_512), .B1 (n_1_687), .B2 (n_1_547), .C1 (n_1_617), .C2 (n_1_572));
OAI22_X1 i_1_702 (.ZN (n_1_510), .A1 (n_1_608), .A2 (n_1_538), .B1 (n_1_681), .B2 (n_1_584));
INV_X1 i_1_701 (.ZN (n_1_509), .A (n_1_510));
OAI221_X1 i_1_700 (.ZN (n_1_508), .A (n_1_509), .B1 (n_1_599), .B2 (n_1_550), .C1 (n_1_652), .C2 (n_1_578));
OAI22_X1 i_1_699 (.ZN (n_1_507), .A1 (n_1_603), .A2 (n_1_531), .B1 (n_1_612), .B2 (n_1_566));
INV_X1 i_1_698 (.ZN (n_1_506), .A (n_1_507));
NOR2_X1 i_1_697 (.ZN (n_1_505), .A1 (n_1_779), .A2 (n_1_663));
INV_X2 i_1_696 (.ZN (n_1_504), .A (n_1_505));
OAI221_X1 i_1_695 (.ZN (n_1_503), .A (n_1_506), .B1 (n_1_656), .B2 (n_1_560), .C1 (n_1_563), .C2 (n_1_504));
OAI22_X1 i_1_694 (.ZN (n_1_502), .A1 (n_1_673), .A2 (n_1_581), .B1 (CLOCK_sgo__n273), .B2 (n_1_553));
INV_X1 i_1_693 (.ZN (n_1_501), .A (n_1_502));
OAI221_X1 i_1_692 (.ZN (n_1_500), .A (n_1_501), .B1 (n_1_621), .B2 (n_1_556), .C1 (n_1_632), .C2 (n_1_541));
OR4_X1 i_1_691 (.ZN (n_1_499), .A1 (n_1_511), .A2 (n_1_508), .A3 (n_1_503), .A4 (n_1_500));
OR3_X1 i_1_690 (.ZN (n_261), .A1 (n_1_718), .A2 (n_1_499), .A3 (n_1_514));
OAI22_X1 i_1_689 (.ZN (n_1_498), .A1 (n_1_664), .A2 (n_1_628), .B1 (n_1_652), .B2 (n_1_600));
INV_X1 i_1_688 (.ZN (n_1_497), .A (n_1_498));
OAI221_X1 i_1_687 (.ZN (n_1_496), .A (n_1_497), .B1 (n_1_674), .B2 (n_1_603), .C1 (n_1_656), .C2 (n_1_637));
AOI22_X1 i_1_686 (.ZN (n_1_495), .A1 (n_1_654), .A2 (n_1_505), .B1 (n_1_633), .B2 (n_1_626));
OAI221_X1 i_1_685 (.ZN (n_1_494), .A (n_1_495), .B1 (n_1_618), .B2 (n_1_617), .C1 (n_1_621), .C2 (n_1_605));
OAI222_X1 i_1_684 (.ZN (n_1_493), .A1 (n_1_684), .A2 (n_1_673), .B1 (n_1_629), .B2 (n_1_599)
    , .C1 (n_1_608), .C2 (n_1_596));
OAI22_X1 i_1_683 (.ZN (n_1_492), .A1 (n_1_678), .A2 (n_1_667), .B1 (CLOCK_sgo__n273), .B2 (n_1_609));
INV_X1 i_1_682 (.ZN (n_1_491), .A (n_1_492));
OAI221_X1 i_1_681 (.ZN (n_1_490), .A (n_1_491), .B1 (n_1_687), .B2 (n_1_649), .C1 (n_1_670), .C2 (n_1_612));
OR4_X1 i_1_680 (.ZN (n_1_489), .A1 (n_1_496), .A2 (n_1_494), .A3 (n_1_493), .A4 (n_1_490));
OR3_X1 i_1_679 (.ZN (n_260), .A1 (n_1_718), .A2 (n_1_489), .A3 (n_1_514));
NOR2_X1 i_1_678 (.ZN (n_1_488), .A1 (n_1_690), .A2 (n_1_587));
NOR2_X2 i_1_677 (.ZN (n_1_487), .A1 (n_1_722), .A2 (n_1_716));
INV_X1 i_1_676 (.ZN (n_1_486), .A (n_1_487));
NOR2_X1 i_1_675 (.ZN (n_1_485), .A1 (n_1_644), .A2 (n_1_487));
OAI21_X1 i_1_674 (.ZN (n_1_484), .A (n_1_488), .B1 (n_1_728), .B2 (n_1_485));
OAI22_X1 i_1_673 (.ZN (n_1_483), .A1 (n_1_687), .A2 (n_1_534), .B1 (n_1_572), .B2 (n_1_504));
INV_X1 i_1_672 (.ZN (n_1_482), .A (n_1_483));
OAI221_X1 i_1_671 (.ZN (n_1_481), .A (n_1_482), .B1 (n_1_632), .B2 (n_1_547), .C1 (CLOCK_sgo__n273), .C2 (n_1_538));
OAI22_X1 i_1_670 (.ZN (n_1_480), .A1 (n_1_667), .A2 (n_1_531), .B1 (n_1_603), .B2 (n_1_584));
INV_X1 i_1_669 (.ZN (n_1_479), .A (n_1_480));
OAI221_X1 i_1_668 (.ZN (n_1_478), .A (n_1_479), .B1 (n_1_617), .B2 (n_1_560), .C1 (n_1_608), .C2 (n_1_566));
OAI22_X1 i_1_667 (.ZN (n_1_477), .A1 (n_1_628), .A2 (n_1_578), .B1 (n_1_599), .B2 (n_1_581));
INV_X1 i_1_666 (.ZN (n_1_476), .A (n_1_477));
OAI221_X1 i_1_665 (.ZN (n_1_475), .A (n_1_476), .B1 (n_1_612), .B2 (n_1_550), .C1 (n_1_673), .C2 (n_1_541));
OAI22_X1 i_1_664 (.ZN (n_1_474), .A1 (n_1_621), .A2 (n_1_553), .B1 (n_1_652), .B2 (n_1_575));
OAI22_X1 i_1_663 (.ZN (n_1_473), .A1 (n_1_656), .A2 (n_1_556), .B1 (n_1_563), .B2 (n_1_516));
OR2_X1 i_1_662 (.ZN (n_1_472), .A1 (n_1_700), .A2 (n_1_593));
OR4_X1 i_1_661 (.ZN (n_1_471), .A1 (n_1_474), .A2 (n_1_473), .A3 (n_1_475), .A4 (n_1_472));
OR4_X1 i_1_660 (.ZN (n_259), .A1 (n_1_481), .A2 (n_1_478), .A3 (n_1_471), .A4 (n_1_484));
OAI22_X1 i_1_659 (.ZN (n_1_470), .A1 (n_1_678), .A2 (n_1_652), .B1 (n_1_653), .B2 (n_1_516));
INV_X1 i_1_658 (.ZN (n_1_469), .A (n_1_470));
OAI221_X1 i_1_657 (.ZN (n_1_468), .A (n_1_469), .B1 (n_1_673), .B2 (n_1_625), .C1 (n_1_670), .C2 (n_1_608));
OAI22_X1 i_1_656 (.ZN (n_1_467), .A1 (n_1_687), .A2 (n_1_664), .B1 (n_1_637), .B2 (n_1_617));
INV_X1 i_1_655 (.ZN (n_1_466), .A (n_1_467));
OAI221_X1 i_1_654 (.ZN (n_1_465), .A (n_1_466), .B1 (n_1_656), .B2 (n_1_605), .C1 (n_1_621), .C2 (n_1_609));
OAI222_X1 i_1_653 (.ZN (n_1_464), .A1 (n_1_628), .A2 (n_1_600), .B1 (CLOCK_sgo__n273)
    , .B2 (n_1_596), .C1 (n_1_684), .C2 (n_1_599));
OAI22_X1 i_1_652 (.ZN (n_1_463), .A1 (n_1_629), .A2 (n_1_612), .B1 (n_1_649), .B2 (n_1_632));
OAI22_X1 i_1_651 (.ZN (n_1_462), .A1 (n_1_674), .A2 (n_1_667), .B1 (n_1_618), .B2 (n_1_504));
OR4_X1 i_1_650 (.ZN (n_1_461), .A1 (n_1_463), .A2 (n_1_462), .A3 (n_1_464), .A4 (n_1_472));
OR4_X1 i_1_649 (.ZN (n_258), .A1 (n_1_468), .A2 (n_1_465), .A3 (n_1_461), .A4 (n_1_484));
OAI222_X1 i_1_648 (.ZN (n_1_460), .A1 (n_1_599), .A2 (n_1_541), .B1 (n_1_608), .B2 (n_1_550)
    , .C1 (n_1_652), .C2 (n_1_531));
NOR3_X1 i_1_647 (.ZN (n_1_459), .A1 (n_1_700), .A2 (n_1_460), .A3 (n_1_593));
OAI22_X1 i_1_646 (.ZN (n_1_458), .A1 (n_1_612), .A2 (n_1_581), .B1 (n_1_687), .B2 (n_1_578));
AOI221_X1 i_1_645 (.ZN (n_1_457), .A (n_1_458), .B1 (n_1_633), .B2 (n_1_535), .C1 (n_1_616), .C2 (n_1_557));
OAI221_X1 i_1_644 (.ZN (n_1_456), .A (n_1_457), .B1 (n_1_560), .B2 (n_1_504), .C1 (n_1_667), .C2 (n_1_584));
OAI21_X1 i_1_643 (.ZN (n_1_455), .A (n_1_729), .B1 (n_1_646), .B2 (n_1_487));
OAI21_X1 i_1_642 (.ZN (n_1_454), .A (n_1_455), .B1 (n_1_572), .B2 (n_1_516));
INV_X1 i_1_641 (.ZN (n_1_453), .A (n_1_454));
OAI221_X1 i_1_640 (.ZN (n_1_452), .A (n_1_453), .B1 (n_1_656), .B2 (n_1_553), .C1 (CLOCK_sgo__n273), .C2 (n_1_566));
OAI22_X1 i_1_639 (.ZN (n_1_451), .A1 (n_1_621), .A2 (n_1_538), .B1 (n_1_647), .B2 (n_1_563));
OAI22_X1 i_1_638 (.ZN (n_1_450), .A1 (n_1_628), .A2 (n_1_575), .B1 (n_1_673), .B2 (n_1_547));
NOR4_X1 i_1_637 (.ZN (n_1_449), .A1 (n_1_451), .A2 (n_1_450), .A3 (n_1_452), .A4 (n_1_456));
NAND3_X1 i_1_636 (.ZN (n_257), .A1 (n_1_488), .A2 (n_1_449), .A3 (n_1_459));
OAI21_X1 i_1_635 (.ZN (n_1_448), .A (n_1_455), .B1 (n_1_625), .B2 (n_1_599));
INV_X1 i_1_634 (.ZN (n_1_447), .A (n_1_448));
OAI221_X1 i_1_633 (.ZN (n_1_446), .A (n_1_447), .B1 (n_1_664), .B2 (n_1_632), .C1 (n_1_687), .C2 (n_1_600));
OAI22_X1 i_1_632 (.ZN (n_1_445), .A1 (n_1_678), .A2 (n_1_628), .B1 (n_1_653), .B2 (n_1_647));
INV_X1 i_1_631 (.ZN (n_1_444), .A (n_1_445));
OAI221_X1 i_1_630 (.ZN (n_1_443), .A (n_1_444), .B1 (n_1_656), .B2 (n_1_609), .C1 (n_1_637), .C2 (n_1_504));
AOI22_X1 i_1_629 (.ZN (n_1_442), .A1 (n_1_616), .A2 (n_1_606), .B1 (n_1_619), .B2 (n_1_517));
OAI221_X1 i_1_628 (.ZN (n_1_441), .A (n_1_442), .B1 (n_1_621), .B2 (n_1_596), .C1 (n_1_674), .C2 (n_1_652));
OAI22_X1 i_1_627 (.ZN (n_1_440), .A1 (n_1_673), .A2 (n_1_649), .B1 (n_1_684), .B2 (n_1_612));
INV_X1 i_1_626 (.ZN (n_1_439), .A (n_1_440));
OAI221_X1 i_1_625 (.ZN (n_1_438), .A (n_1_439), .B1 (n_1_629), .B2 (n_1_608), .C1 (n_1_670), .C2 (n_1_640));
OR4_X1 i_1_624 (.ZN (n_1_437), .A1 (n_1_443), .A2 (n_1_441), .A3 (n_1_586), .A4 (n_1_438));
OR4_X1 i_1_623 (.ZN (n_256), .A1 (n_1_705), .A2 (n_1_446), .A3 (n_1_437), .A4 (n_1_591));
OAI22_X1 i_1_622 (.ZN (n_1_436), .A1 (n_1_621), .A2 (n_1_566), .B1 (n_1_673), .B2 (n_1_534));
OAI22_X1 i_1_621 (.ZN (n_1_435), .A1 (n_1_632), .A2 (n_1_578), .B1 (n_1_645), .B2 (n_1_563));
OAI22_X1 i_1_620 (.ZN (n_1_434), .A1 (n_1_617), .A2 (n_1_553), .B1 (n_1_652), .B2 (n_1_584));
OAI22_X1 i_1_619 (.ZN (n_1_433), .A1 (n_1_628), .A2 (n_1_531), .B1 (n_1_556), .B2 (n_1_504));
OR4_X1 i_1_618 (.ZN (n_1_432), .A1 (n_1_436), .A2 (n_1_435), .A3 (n_1_434), .A4 (n_1_433));
OAI22_X1 i_1_617 (.ZN (n_1_431), .A1 (n_1_599), .A2 (n_1_547), .B1 (n_1_612), .B2 (n_1_541));
INV_X1 i_1_616 (.ZN (n_1_430), .A (n_1_431));
OAI221_X1 i_1_615 (.ZN (n_1_429), .A (n_1_430), .B1 (n_1_608), .B2 (n_1_581), .C1 (n_1_560), .C2 (n_1_516));
OAI22_X1 i_1_614 (.ZN (n_1_428), .A1 (n_1_687), .A2 (n_1_575), .B1 (n_1_656), .B2 (n_1_538));
INV_X1 i_1_613 (.ZN (n_1_427), .A (n_1_428));
OAI221_X1 i_1_612 (.ZN (n_1_426), .A (n_1_427), .B1 (n_1_647), .B2 (n_1_572), .C1 (CLOCK_sgo__n273), .C2 (n_1_550));
OR4_X1 i_1_611 (.ZN (n_255), .A1 (n_1_429), .A2 (n_1_426), .A3 (n_1_432), .A4 (n_1_585));
OAI22_X1 i_1_610 (.ZN (n_1_425), .A1 (n_1_670), .A2 (n_1_621), .B1 (n_1_673), .B2 (n_1_664));
OAI22_X1 i_1_609 (.ZN (n_1_424), .A1 (CLOCK_sgo__n273), .A2 (n_1_629), .B1 (n_1_674), .B2 (n_1_628));
OR4_X1 i_1_608 (.ZN (n_1_423), .A1 (n_1_425), .A2 (n_1_424), .A3 (n_1_590), .A4 (n_1_587));
OAI22_X1 i_1_607 (.ZN (n_1_422), .A1 (n_1_653), .A2 (n_1_645), .B1 (n_1_649), .B2 (n_1_599));
INV_X1 i_1_606 (.ZN (n_1_421), .A (n_1_422));
OAI221_X1 i_1_605 (.ZN (n_1_420), .A (n_1_421), .B1 (n_1_647), .B2 (n_1_618), .C1 (n_1_625), .C2 (n_1_612));
AOI22_X1 i_1_604 (.ZN (n_1_419), .A1 (n_1_616), .A2 (n_1_610), .B1 (n_1_633), .B2 (n_1_601));
OAI221_X1 i_1_603 (.ZN (n_1_418), .A (n_1_419), .B1 (n_1_656), .B2 (n_1_596), .C1 (n_1_605), .C2 (n_1_504));
OAI222_X1 i_1_602 (.ZN (n_1_417), .A1 (n_1_637), .A2 (n_1_516), .B1 (n_1_687), .B2 (n_1_678)
    , .C1 (n_1_684), .C2 (n_1_608));
OR4_X1 i_1_601 (.ZN (n_1_416), .A1 (n_1_420), .A2 (n_1_418), .A3 (n_1_700), .A4 (n_1_417));
OR3_X1 i_1_600 (.ZN (n_254), .A1 (n_1_423), .A2 (n_1_416), .A3 (n_1_591));
OAI22_X1 i_1_599 (.ZN (n_1_415), .A1 (n_1_661), .A2 (n_1_563), .B1 (n_1_556), .B2 (n_1_516));
OAI22_X1 i_1_598 (.ZN (n_1_414), .A1 (n_1_621), .A2 (n_1_550), .B1 (n_1_647), .B2 (n_1_560));
OAI22_X1 i_1_597 (.ZN (n_1_413), .A1 (n_1_687), .A2 (n_1_531), .B1 (n_1_628), .B2 (n_1_584));
OAI22_X1 i_1_596 (.ZN (n_1_412), .A1 (n_1_673), .A2 (n_1_578), .B1 (n_1_553), .B2 (n_1_504));
OR4_X1 i_1_595 (.ZN (n_1_411), .A1 (n_1_415), .A2 (n_1_414), .A3 (n_1_413), .A4 (n_1_412));
OAI22_X1 i_1_594 (.ZN (n_1_410), .A1 (n_1_608), .A2 (n_1_541), .B1 (n_1_656), .B2 (n_1_566));
INV_X1 i_1_593 (.ZN (n_1_409), .A (n_1_410));
OAI221_X1 i_1_592 (.ZN (n_1_408), .A (n_1_409), .B1 (n_1_612), .B2 (n_1_547), .C1 (n_1_617), .C2 (n_1_538));
AOI22_X1 i_1_591 (.ZN (n_1_407), .A1 (n_1_633), .A2 (n_1_576), .B1 (n_1_646), .B2 (n_1_573));
OAI221_X1 i_1_590 (.ZN (n_1_406), .A (n_1_407), .B1 (n_1_599), .B2 (n_1_534), .C1 (CLOCK_sgo__n273), .C2 (n_1_581));
OR4_X1 i_1_589 (.ZN (n_253), .A1 (n_1_408), .A2 (n_1_406), .A3 (n_1_411), .A4 (n_1_688));
OAI222_X1 i_1_588 (.ZN (n_1_405), .A1 (n_1_661), .A2 (n_1_653), .B1 (n_1_678), .B2 (n_1_632)
    , .C1 (n_1_625), .C2 (n_1_608));
OR3_X1 i_1_587 (.ZN (n_1_404), .A1 (n_1_711), .A2 (n_1_938), .A3 (n_1_590));
OAI22_X1 i_1_586 (.ZN (n_1_403), .A1 (n_1_647), .A2 (n_1_637), .B1 (n_1_649), .B2 (n_1_612));
OAI22_X1 i_1_585 (.ZN (n_1_402), .A1 (n_1_645), .A2 (n_1_618), .B1 (n_1_664), .B2 (n_1_599));
OR4_X1 i_1_584 (.ZN (n_1_401), .A1 (n_1_723), .A2 (n_1_706), .A3 (n_1_403), .A4 (n_1_402));
OAI22_X1 i_1_583 (.ZN (n_1_400), .A1 (n_1_609), .A2 (n_1_504), .B1 (n_1_673), .B2 (n_1_600));
INV_X1 i_1_582 (.ZN (n_1_399), .A (n_1_400));
OAI221_X1 i_1_581 (.ZN (n_1_398), .A (n_1_399), .B1 (n_1_629), .B2 (n_1_621), .C1 (n_1_617), .C2 (n_1_596));
OAI22_X1 i_1_580 (.ZN (n_1_397), .A1 (n_1_687), .A2 (n_1_674), .B1 (n_1_670), .B2 (n_1_656));
INV_X1 i_1_579 (.ZN (n_1_396), .A (n_1_397));
OAI221_X1 i_1_578 (.ZN (n_1_395), .A (n_1_396), .B1 (n_1_684), .B2 (n_1_640), .C1 (n_1_605), .C2 (n_1_516));
OR4_X1 i_1_577 (.ZN (n_1_394), .A1 (n_1_398), .A2 (n_1_395), .A3 (n_1_401), .A4 (n_1_404));
OR4_X1 i_1_576 (.ZN (n_252), .A1 (n_1_690), .A2 (n_1_405), .A3 (n_1_593), .A4 (n_1_394));
OR2_X1 i_1_575 (.ZN (n_1_393), .A1 (n_1_691), .A2 (n_1_593));
OR2_X1 i_1_574 (.ZN (n_1_392), .A1 (n_1_706), .A2 (n_1_393));
OAI22_X1 i_1_573 (.ZN (n_1_391), .A1 (n_1_612), .A2 (n_1_534), .B1 (n_1_724), .B2 (n_1_563));
INV_X1 i_1_572 (.ZN (n_1_390), .A (n_1_391));
OAI221_X1 i_1_571 (.ZN (n_1_389), .A (n_1_390), .B1 (n_1_538), .B2 (n_1_504), .C1 (n_1_617), .C2 (n_1_566));
OAI22_X1 i_1_570 (.ZN (n_1_388), .A1 (n_1_656), .A2 (n_1_550), .B1 (n_1_673), .B2 (n_1_575));
INV_X1 i_1_569 (.ZN (n_1_387), .A (n_1_388));
OAI221_X1 i_1_568 (.ZN (n_1_386), .A (n_1_387), .B1 (n_1_621), .B2 (n_1_581), .C1 (n_1_608), .C2 (n_1_547));
OAI22_X1 i_1_567 (.ZN (n_1_385), .A1 (n_1_647), .A2 (n_1_556), .B1 (n_1_632), .B2 (n_1_531));
OAI22_X1 i_1_566 (.ZN (n_1_384), .A1 (n_1_599), .A2 (n_1_578), .B1 (n_1_553), .B2 (n_1_516));
OR4_X1 i_1_565 (.ZN (n_1_383), .A1 (n_1_385), .A2 (n_1_384), .A3 (n_1_386), .A4 (n_1_389));
AOI22_X1 i_1_564 (.ZN (n_1_382), .A1 (n_1_662), .A2 (n_1_573), .B1 (n_1_646), .B2 (n_1_561));
OAI221_X1 i_1_563 (.ZN (n_1_381), .A (n_1_382), .B1 (n_1_640), .B2 (n_1_541), .C1 (n_1_687), .C2 (n_1_584));
OR3_X1 i_1_562 (.ZN (n_1_380), .A1 (n_1_693), .A2 (n_1_381), .A3 (n_1_404));
OR3_X1 i_1_561 (.ZN (n_251), .A1 (n_1_383), .A2 (n_1_380), .A3 (n_1_392));
OAI222_X1 i_1_560 (.ZN (n_1_379), .A1 (n_1_664), .A2 (n_1_612), .B1 (n_1_645), .B2 (n_1_637)
    , .C1 (n_1_661), .C2 (n_1_618));
OAI22_X1 i_1_559 (.ZN (n_1_378), .A1 (n_1_600), .A2 (n_1_599), .B1 (n_1_647), .B2 (n_1_605));
OAI22_X1 i_1_558 (.ZN (n_1_377), .A1 (n_1_684), .A2 (n_1_621), .B1 (n_1_649), .B2 (n_1_608));
NOR4_X1 i_1_557 (.ZN (n_1_376), .A1 (n_1_378), .A2 (n_1_377), .A3 (n_1_379), .A4 (n_1_719));
OAI22_X1 i_1_556 (.ZN (n_1_375), .A1 (n_1_640), .A2 (n_1_625), .B1 (n_1_609), .B2 (n_1_516));
OAI22_X1 i_1_555 (.ZN (n_1_374), .A1 (n_1_678), .A2 (n_1_673), .B1 (n_1_596), .B2 (n_1_504));
OAI22_X1 i_1_554 (.ZN (n_1_373), .A1 (n_1_670), .A2 (n_1_617), .B1 (n_1_724), .B2 (n_1_653));
OAI22_X1 i_1_553 (.ZN (n_1_372), .A1 (n_1_674), .A2 (n_1_632), .B1 (n_1_656), .B2 (n_1_629));
NOR4_X1 i_1_552 (.ZN (n_1_371), .A1 (n_1_375), .A2 (n_1_374), .A3 (n_1_373), .A4 (n_1_372));
NAND3_X1 i_1_551 (.ZN (n_250), .A1 (n_1_689), .A2 (n_1_371), .A3 (n_1_376));
OR3_X1 i_1_550 (.ZN (n_1_370), .A1 (n_1_703), .A2 (n_1_690), .A3 (n_1_589));
OAI22_X1 i_1_549 (.ZN (n_1_369), .A1 (n_1_566), .A2 (n_1_504), .B1 (n_1_673), .B2 (n_1_531));
INV_X1 i_1_548 (.ZN (n_1_368), .A (n_1_369));
OAI221_X1 i_1_547 (.ZN (n_1_367), .A (n_1_368), .B1 (n_1_617), .B2 (n_1_550), .C1 (n_1_621), .C2 (n_1_541));
OAI22_X1 i_1_546 (.ZN (n_1_366), .A1 (n_1_647), .A2 (n_1_553), .B1 (n_1_632), .B2 (n_1_584));
INV_X1 i_1_545 (.ZN (n_1_365), .A (n_1_366));
OAI221_X1 i_1_544 (.ZN (n_1_364), .A (n_1_365), .B1 (n_1_724), .B2 (n_1_572), .C1 (n_1_608), .C2 (n_1_534));
AOI22_X1 i_1_543 (.ZN (n_1_363), .A1 (n_1_662), .A2 (n_1_561), .B1 (n_1_646), .B2 (n_1_557));
OAI221_X1 i_1_542 (.ZN (n_1_362), .A (n_1_363), .B1 (n_1_701), .B2 (n_1_563), .C1 (n_1_656), .C2 (n_1_581));
OAI22_X1 i_1_541 (.ZN (n_1_361), .A1 (n_1_538), .A2 (n_1_516), .B1 (n_1_640), .B2 (n_1_547));
OAI22_X1 i_1_540 (.ZN (n_1_360), .A1 (n_1_599), .A2 (n_1_575), .B1 (n_1_612), .B2 (n_1_578));
OR4_X1 i_1_539 (.ZN (n_1_359), .A1 (n_1_361), .A2 (n_1_360), .A3 (n_1_362), .A4 (n_1_593));
OR4_X1 i_1_538 (.ZN (n_249), .A1 (n_1_367), .A2 (n_1_364), .A3 (n_1_359), .A4 (n_1_370));
OAI22_X1 i_1_537 (.ZN (n_1_358), .A1 (n_1_701), .A2 (n_1_653), .B1 (n_1_678), .B2 (n_1_599));
INV_X1 i_1_536 (.ZN (n_1_357), .A (n_1_358));
OAI221_X1 i_1_535 (.ZN (n_1_356), .A (n_1_357), .B1 (n_1_661), .B2 (n_1_637), .C1 (n_1_724), .C2 (n_1_618));
OAI22_X1 i_1_534 (.ZN (n_1_355), .A1 (n_1_649), .A2 (n_1_640), .B1 (n_1_645), .B2 (n_1_605));
INV_X1 i_1_533 (.ZN (n_1_354), .A (n_1_355));
OAI221_X1 i_1_532 (.ZN (n_1_353), .A (n_1_354), .B1 (n_1_684), .B2 (n_1_656), .C1 (n_1_664), .C2 (n_1_608));
OAI222_X1 i_1_531 (.ZN (n_1_352), .A1 (n_1_612), .A2 (n_1_600), .B1 (n_1_674), .B2 (n_1_673)
    , .C1 (n_1_647), .C2 (n_1_609));
OAI22_X1 i_1_530 (.ZN (n_1_351), .A1 (n_1_596), .A2 (n_1_516), .B1 (n_1_670), .B2 (n_1_504));
OAI22_X1 i_1_529 (.ZN (n_1_350), .A1 (n_1_629), .A2 (n_1_617), .B1 (n_1_625), .B2 (n_1_621));
OR4_X1 i_1_528 (.ZN (n_1_349), .A1 (n_1_351), .A2 (n_1_350), .A3 (n_1_352), .A4 (n_1_593));
OR4_X1 i_1_527 (.ZN (n_248), .A1 (n_1_356), .A2 (n_1_353), .A3 (n_1_349), .A4 (n_1_370));
OAI22_X1 i_1_526 (.ZN (n_1_348), .A1 (CLOCK_sgo__n273), .A2 (n_1_534), .B1 (n_1_647), .B2 (n_1_538));
OAI22_X1 i_1_525 (.ZN (n_1_347), .A1 (n_1_656), .A2 (n_1_541), .B1 (n_1_617), .B2 (n_1_581));
OAI22_X1 i_1_524 (.ZN (n_1_346), .A1 (n_1_599), .A2 (n_1_531), .B1 (n_1_673), .B2 (n_1_584));
OAI22_X1 i_1_523 (.ZN (n_1_345), .A1 (n_1_724), .A2 (n_1_560), .B1 (n_1_621), .B2 (n_1_547));
OR4_X1 i_1_522 (.ZN (n_1_344), .A1 (n_1_348), .A2 (n_1_347), .A3 (n_1_346), .A4 (n_1_345));
AOI22_X1 i_1_521 (.ZN (n_1_343), .A1 (n_1_646), .A2 (n_1_554), .B1 (n_1_567), .B2 (n_1_517));
OAI221_X1 i_1_520 (.ZN (n_1_342), .A (n_1_343), .B1 (n_1_608), .B2 (n_1_578), .C1 (n_1_550), .C2 (n_1_504));
OAI22_X1 i_1_519 (.ZN (n_1_341), .A1 (n_1_701), .A2 (n_1_572), .B1 (n_1_704), .B2 (n_1_563));
INV_X1 i_1_518 (.ZN (n_1_340), .A (n_1_341));
OAI221_X1 i_1_517 (.ZN (n_1_339), .A (n_1_340), .B1 (n_1_612), .B2 (n_1_575), .C1 (n_1_661), .C2 (n_1_556));
OR4_X1 i_1_516 (.ZN (n_247), .A1 (n_1_342), .A2 (n_1_339), .A3 (n_1_344), .A4 (n_1_588));
AOI22_X1 i_1_515 (.ZN (n_1_338), .A1 (n_1_662), .A2 (n_1_606), .B1 (n_1_646), .B2 (n_1_610));
OAI221_X1 i_1_514 (.ZN (n_1_337), .A (n_1_338), .B1 (n_1_629), .B2 (n_1_504), .C1 (n_1_684), .C2 (n_1_617));
AOI22_X1 i_1_513 (.ZN (n_1_336), .A1 (n_1_725), .A2 (n_1_638), .B1 (n_1_650), .B2 (n_1_622));
OAI221_X1 i_1_512 (.ZN (n_1_335), .A (n_1_336), .B1 (n_1_656), .B2 (n_1_625), .C1 (n_1_670), .C2 (n_1_516));
NOR2_X1 i_1_511 (.ZN (n_1_334), .A1 (n_1_674), .A2 (n_1_599));
OAI22_X1 i_1_510 (.ZN (n_1_333), .A1 (n_1_701), .A2 (n_1_618), .B1 (n_1_664), .B2 (n_1_640));
OAI22_X1 i_1_509 (.ZN (n_1_332), .A1 (n_1_678), .A2 (n_1_612), .B1 (n_1_608), .B2 (n_1_600));
OAI22_X1 i_1_508 (.ZN (n_1_331), .A1 (n_1_704), .A2 (n_1_653), .B1 (n_1_647), .B2 (n_1_596));
OR4_X1 i_1_507 (.ZN (n_1_330), .A1 (n_1_334), .A2 (n_1_333), .A3 (n_1_332), .A4 (n_1_331));
OR4_X1 i_1_506 (.ZN (n_246), .A1 (n_1_337), .A2 (n_1_335), .A3 (n_1_330), .A4 (n_1_588));
OAI22_X1 i_1_505 (.ZN (n_1_329), .A1 (n_1_608), .A2 (n_1_575), .B1 (n_1_599), .B2 (n_1_584));
INV_X1 i_1_504 (.ZN (n_1_328), .A (n_1_329));
OAI221_X1 i_1_503 (.ZN (n_1_327), .A (n_1_328), .B1 (n_1_581), .B2 (n_1_504), .C1 (n_1_724), .C2 (n_1_556));
AOI22_X1 i_1_502 (.ZN (n_1_326), .A1 (n_1_662), .A2 (n_1_554), .B1 (n_1_564), .B2 (n_1_487));
OAI221_X1 i_1_501 (.ZN (n_1_325), .A (n_1_326), .B1 (n_1_550), .B2 (n_1_516), .C1 (n_1_656), .C2 (n_1_547));
OAI22_X1 i_1_500 (.ZN (n_1_324), .A1 (n_1_617), .A2 (n_1_541), .B1 (n_1_701), .B2 (n_1_560));
OAI22_X1 i_1_499 (.ZN (n_1_323), .A1 (n_1_612), .A2 (n_1_531), .B1 (n_1_621), .B2 (n_1_534));
AOI22_X1 i_1_498 (.ZN (n_1_322), .A1 (n_1_646), .A2 (n_1_539), .B1 (n_1_648), .B2 (n_1_567));
OAI221_X1 i_1_497 (.ZN (n_1_321), .A (n_1_322), .B1 (n_1_640), .B2 (n_1_578), .C1 (n_1_704), .C2 (n_1_572));
OR4_X1 i_1_496 (.ZN (n_1_320), .A1 (n_1_324), .A2 (n_1_323), .A3 (n_1_321), .A4 (n_1_325));
OR4_X1 i_1_495 (.ZN (n_245), .A1 (n_1_705), .A2 (n_1_327), .A3 (n_1_320), .A4 (n_1_591));
OAI21_X1 i_1_494 (.ZN (n_1_319), .A (n_1_710), .B1 (n_1_656), .B2 (n_1_649));
INV_X1 i_1_493 (.ZN (n_1_318), .A (n_1_319));
OAI221_X1 i_1_492 (.ZN (n_1_317), .A (n_1_318), .B1 (n_1_640), .B2 (n_1_600), .C1 (n_1_664), .C2 (n_1_621));
AOI22_X1 i_1_491 (.ZN (n_1_316), .A1 (n_1_662), .A2 (n_1_610), .B1 (n_1_630), .B2 (n_1_517));
OAI221_X1 i_1_490 (.ZN (n_1_315), .A (n_1_316), .B1 (n_1_724), .B2 (n_1_605), .C1 (n_1_625), .C2 (n_1_617));
OAI22_X1 i_1_489 (.ZN (n_1_314), .A1 (n_1_678), .A2 (n_1_608), .B1 (n_1_704), .B2 (n_1_618));
INV_X1 i_1_488 (.ZN (n_1_313), .A (n_1_314));
OAI221_X1 i_1_487 (.ZN (n_1_312), .A (n_1_313), .B1 (n_1_684), .B2 (n_1_504), .C1 (n_1_701), .C2 (n_1_637));
OAI22_X1 i_1_486 (.ZN (n_1_311), .A1 (n_1_645), .A2 (n_1_596), .B1 (n_1_670), .B2 (n_1_647));
OAI22_X1 i_1_485 (.ZN (n_1_310), .A1 (n_1_653), .A2 (n_1_486), .B1 (n_1_674), .B2 (n_1_612));
OR4_X1 i_1_484 (.ZN (n_1_309), .A1 (n_1_311), .A2 (n_1_310), .A3 (n_1_312), .A4 (n_1_315));
OR4_X1 i_1_483 (.ZN (n_244), .A1 (n_1_693), .A2 (n_1_317), .A3 (n_1_309), .A4 (n_1_392));
OAI22_X1 i_1_482 (.ZN (n_1_308), .A1 (n_1_608), .A2 (n_1_531), .B1 (n_1_645), .B2 (n_1_566));
INV_X1 i_1_481 (.ZN (n_1_307), .A (n_1_308));
OAI221_X1 i_1_480 (.ZN (n_1_306), .A (n_1_307), .B1 (n_1_617), .B2 (n_1_547), .C1 (n_1_612), .C2 (n_1_584));
AOI22_X1 i_1_479 (.ZN (n_1_305), .A1 (n_1_542), .A2 (n_1_505), .B1 (n_1_712), .B2 (n_1_564));
OAI221_X1 i_1_478 (.ZN (n_1_304), .A (n_1_305), .B1 (n_1_661), .B2 (n_1_538), .C1 (n_1_724), .C2 (n_1_553));
AOI22_X1 i_1_477 (.ZN (n_1_303), .A1 (n_1_582), .A2 (n_1_517), .B1 (n_1_573), .B2 (n_1_487));
OAI221_X1 i_1_476 (.ZN (n_1_302), .A (n_1_303), .B1 (n_1_621), .B2 (n_1_578), .C1 (n_1_704), .C2 (n_1_560));
OAI22_X1 i_1_475 (.ZN (n_1_301), .A1 (n_1_656), .A2 (n_1_534), .B1 (n_1_701), .B2 (n_1_556));
OAI22_X1 i_1_474 (.ZN (n_1_300), .A1 (n_1_640), .A2 (n_1_575), .B1 (n_1_647), .B2 (n_1_550));
OR4_X1 i_1_473 (.ZN (n_1_299), .A1 (n_1_301), .A2 (n_1_300), .A3 (n_1_302), .A4 (n_1_304));
OR4_X1 i_1_472 (.ZN (n_243), .A1 (n_1_693), .A2 (n_1_306), .A3 (n_1_299), .A4 (n_1_392));
OR2_X1 i_1_471 (.ZN (n_1_298), .A1 (n_1_695), .A2 (n_1_393));
OAI22_X1 i_1_470 (.ZN (n_1_297), .A1 (n_1_647), .A2 (n_1_629), .B1 (n_1_621), .B2 (n_1_600));
OAI22_X1 i_1_469 (.ZN (n_1_296), .A1 (n_1_713), .A2 (n_1_653), .B1 (n_1_649), .B2 (n_1_617));
OR4_X1 i_1_468 (.ZN (n_1_295), .A1 (n_1_706), .A2 (n_1_699), .A3 (n_1_297), .A4 (n_1_296));
OAI222_X1 i_1_467 (.ZN (n_1_294), .A1 (n_1_661), .A2 (n_1_596), .B1 (n_1_625), .B2 (n_1_504)
    , .C1 (n_1_724), .C2 (n_1_609));
OAI22_X1 i_1_466 (.ZN (n_1_293), .A1 (n_1_678), .A2 (n_1_640), .B1 (n_1_670), .B2 (n_1_645));
INV_X1 i_1_465 (.ZN (n_1_292), .A (n_1_293));
OAI221_X1 i_1_464 (.ZN (n_1_291), .A (n_1_292), .B1 (n_1_664), .B2 (n_1_656), .C1 (n_1_674), .C2 (n_1_608));
OAI22_X1 i_1_463 (.ZN (n_1_290), .A1 (n_1_684), .A2 (n_1_516), .B1 (n_1_701), .B2 (n_1_605));
OAI22_X1 i_1_462 (.ZN (n_1_289), .A1 (n_1_618), .A2 (n_1_486), .B1 (n_1_704), .B2 (n_1_637));
OR4_X1 i_1_461 (.ZN (n_1_288), .A1 (n_1_290), .A2 (n_1_289), .A3 (n_1_291), .A4 (n_1_294));
OR3_X1 i_1_460 (.ZN (n_242), .A1 (n_1_295), .A2 (n_1_288), .A3 (n_1_298));
OAI22_X1 i_1_459 (.ZN (n_1_287), .A1 (n_1_704), .A2 (n_1_556), .B1 (n_1_645), .B2 (n_1_550));
AOI221_X1 i_1_458 (.ZN (n_1_286), .A (n_1_287), .B1 (n_1_622), .B2 (n_1_576), .C1 (n_1_648), .C2 (n_1_582));
OAI211_X1 i_1_457 (.ZN (n_1_285), .A (n_1_698), .B (n_1_286), .C1 (n_1_608), .C2 (n_1_584));
OAI222_X1 i_1_456 (.ZN (n_1_284), .A1 (n_1_724), .A2 (n_1_538), .B1 (n_1_617), .B2 (n_1_534)
    , .C1 (n_1_547), .C2 (n_1_504));
OAI22_X1 i_1_455 (.ZN (n_1_283), .A1 (n_1_560), .A2 (n_1_486), .B1 (CLOCK_sgo__n273), .B2 (n_1_531));
INV_X1 i_1_454 (.ZN (n_1_282), .A (n_1_283));
OAI221_X1 i_1_453 (.ZN (n_1_281), .A (n_1_282), .B1 (n_1_656), .B2 (n_1_578), .C1 (n_1_701), .C2 (n_1_553));
OAI22_X1 i_1_452 (.ZN (n_1_280), .A1 (n_1_541), .A2 (n_1_516), .B1 (n_1_707), .B2 (n_1_563));
OAI22_X1 i_1_451 (.ZN (n_1_279), .A1 (n_1_713), .A2 (n_1_572), .B1 (n_1_661), .B2 (n_1_566));
OR4_X1 i_1_450 (.ZN (n_1_278), .A1 (n_1_280), .A2 (n_1_279), .A3 (n_1_281), .A4 (n_1_284));
OR3_X1 i_1_449 (.ZN (n_241), .A1 (n_1_285), .A2 (n_1_278), .A3 (n_1_298));
AOI22_X1 i_1_448 (.ZN (n_1_277), .A1 (n_1_685), .A2 (n_1_648), .B1 (n_1_708), .B2 (n_1_654));
OAI221_X1 i_1_447 (.ZN (n_1_276), .A (n_1_277), .B1 (n_1_670), .B2 (n_1_661), .C1 (n_1_625), .C2 (n_1_516));
AOI22_X1 i_1_446 (.ZN (n_1_275), .A1 (n_1_725), .A2 (n_1_597), .B1 (n_1_638), .B2 (n_1_487));
OAI221_X1 i_1_445 (.ZN (n_1_274), .A (n_1_275), .B1 (n_1_664), .B2 (n_1_617), .C1 (n_1_713), .C2 (n_1_618));
NOR2_X1 i_1_444 (.ZN (n_1_273), .A1 (n_1_645), .A2 (n_1_629));
OAI22_X1 i_1_443 (.ZN (n_1_272), .A1 (n_1_649), .A2 (n_1_504), .B1 (n_1_656), .B2 (n_1_600));
OAI22_X1 i_1_442 (.ZN (n_1_271), .A1 (n_1_678), .A2 (n_1_621), .B1 (n_1_704), .B2 (n_1_605));
OAI22_X1 i_1_441 (.ZN (n_1_270), .A1 (n_1_674), .A2 (n_1_640), .B1 (n_1_701), .B2 (n_1_609));
OR4_X1 i_1_440 (.ZN (n_1_269), .A1 (n_1_273), .A2 (n_1_272), .A3 (n_1_271), .A4 (n_1_270));
OR4_X1 i_1_439 (.ZN (n_240), .A1 (n_1_276), .A2 (n_1_274), .A3 (n_1_269), .A4 (n_1_591));
OAI22_X1 i_1_438 (.ZN (n_1_268), .A1 (n_1_724), .A2 (n_1_566), .B1 (n_1_534), .B2 (n_1_504));
OAI22_X1 i_1_437 (.ZN (n_1_267), .A1 (n_1_656), .A2 (n_1_575), .B1 (n_1_617), .B2 (n_1_578));
OAI22_X1 i_1_436 (.ZN (n_1_266), .A1 (n_1_547), .A2 (n_1_516), .B1 (n_1_640), .B2 (n_1_584));
OAI22_X1 i_1_435 (.ZN (n_1_265), .A1 (n_1_704), .A2 (n_1_553), .B1 (n_1_661), .B2 (n_1_550));
OR4_X1 i_1_434 (.ZN (n_1_264), .A1 (n_1_268), .A2 (n_1_267), .A3 (n_1_266), .A4 (n_1_265));
AOI22_X1 i_1_433 (.ZN (n_1_263), .A1 (n_1_712), .A2 (n_1_561), .B1 (n_1_708), .B2 (n_1_573));
OAI221_X1 i_1_432 (.ZN (n_1_262), .A (n_1_263), .B1 (n_1_645), .B2 (n_1_581), .C1 (n_1_556), .C2 (n_1_486));
AOI22_X1 i_1_431 (.ZN (n_1_261), .A1 (n_1_648), .A2 (n_1_542), .B1 (n_1_622), .B2 (n_1_532));
OAI221_X1 i_1_430 (.ZN (n_1_260), .A (n_1_261), .B1 (n_1_692), .B2 (n_1_563), .C1 (n_1_701), .C2 (n_1_538));
OR4_X1 i_1_429 (.ZN (n_239), .A1 (n_1_262), .A2 (n_1_260), .A3 (n_1_264), .A4 (n_1_592));
OAI22_X1 i_1_428 (.ZN (n_1_259), .A1 (n_1_684), .A2 (n_1_645), .B1 (n_1_692), .B2 (n_1_653));
INV_X1 i_1_427 (.ZN (n_1_258), .A (n_1_259));
OAI221_X1 i_1_426 (.ZN (n_1_257), .A (n_1_258), .B1 (n_1_605), .B2 (n_1_486), .C1 (n_1_661), .C2 (n_1_629));
OAI22_X1 i_1_425 (.ZN (n_1_256), .A1 (n_1_704), .A2 (n_1_609), .B1 (n_1_713), .B2 (n_1_637));
INV_X1 i_1_424 (.ZN (n_1_255), .A (n_1_256));
OAI221_X1 i_1_423 (.ZN (n_1_254), .A (n_1_255), .B1 (n_1_617), .B2 (n_1_600), .C1 (n_1_674), .C2 (n_1_621));
NOR2_X1 i_1_422 (.ZN (n_1_253), .A1 (n_1_649), .A2 (n_1_516));
OAI22_X1 i_1_421 (.ZN (n_1_252), .A1 (n_1_678), .A2 (n_1_656), .B1 (n_1_707), .B2 (n_1_618));
OAI22_X1 i_1_420 (.ZN (n_1_251), .A1 (n_1_724), .A2 (n_1_670), .B1 (n_1_647), .B2 (n_1_625));
OAI22_X1 i_1_419 (.ZN (n_1_250), .A1 (n_1_701), .A2 (n_1_596), .B1 (n_1_664), .B2 (n_1_504));
OR4_X1 i_1_418 (.ZN (n_1_249), .A1 (n_1_253), .A2 (n_1_252), .A3 (n_1_251), .A4 (n_1_250));
OR4_X1 i_1_417 (.ZN (n_238), .A1 (n_1_257), .A2 (n_1_254), .A3 (n_1_249), .A4 (n_1_592));
NOR3_X4 i_1_416 (.ZN (n_1_248), .A1 (\counter[2] ), .A2 (n_1_717), .A3 (n_1_722));
INV_X1 i_1_415 (.ZN (n_1_247), .A (n_1_248));
AOI22_X1 i_1_414 (.ZN (n_1_246), .A1 (n_1_662), .A2 (n_1_582), .B1 (n_1_554), .B2 (n_1_487));
OAI221_X1 i_1_413 (.ZN (n_1_245), .A (n_1_246), .B1 (n_1_692), .B2 (n_1_572), .C1 (n_1_563), .C2 (n_1_247));
OAI22_X1 i_1_412 (.ZN (n_1_244), .A1 (n_1_713), .A2 (n_1_556), .B1 (n_1_621), .B2 (n_1_584));
OAI22_X1 i_1_411 (.ZN (n_1_243), .A1 (n_1_707), .A2 (n_1_560), .B1 (n_1_645), .B2 (n_1_541));
OAI21_X1 i_1_410 (.ZN (n_1_242), .A (n_1_694), .B1 (n_1_727), .B2 (n_1_721));
AOI22_X1 i_1_409 (.ZN (n_1_241), .A1 (n_1_725), .A2 (n_1_551), .B1 (n_1_648), .B2 (n_1_548));
OAI221_X1 i_1_408 (.ZN (n_1_240), .A (n_1_241), .B1 (n_1_704), .B2 (n_1_538), .C1 (n_1_617), .C2 (n_1_575));
OAI22_X1 i_1_407 (.ZN (n_1_239), .A1 (n_1_578), .A2 (n_1_504), .B1 (n_1_701), .B2 (n_1_566));
OAI22_X1 i_1_406 (.ZN (n_1_238), .A1 (n_1_534), .A2 (n_1_516), .B1 (n_1_656), .B2 (n_1_531));
OR4_X1 i_1_405 (.ZN (n_1_237), .A1 (n_1_239), .A2 (n_1_238), .A3 (n_1_240), .A4 (n_1_242));
OR4_X1 i_1_404 (.ZN (n_237), .A1 (n_1_244), .A2 (n_1_243), .A3 (n_1_245), .A4 (n_1_237));
OAI22_X1 i_1_403 (.ZN (n_1_236), .A1 (n_1_704), .A2 (n_1_596), .B1 (n_1_713), .B2 (n_1_605));
INV_X1 i_1_402 (.ZN (n_1_235), .A (n_1_236));
OAI221_X1 i_1_401 (.ZN (n_1_234), .A (n_1_235), .B1 (n_1_664), .B2 (n_1_516), .C1 (n_1_724), .C2 (n_1_629));
AOI22_X1 i_1_400 (.ZN (n_1_233), .A1 (n_1_679), .A2 (n_1_616), .B1 (n_1_654), .B2 (n_1_248));
OAI221_X1 i_1_399 (.ZN (n_1_232), .A (n_1_233), .B1 (n_1_674), .B2 (n_1_656), .C1 (n_1_701), .C2 (n_1_670));
AOI22_X1 i_1_398 (.ZN (n_1_231), .A1 (n_1_646), .A2 (n_1_626), .B1 (n_1_685), .B2 (n_1_662));
OAI22_X1 i_1_397 (.ZN (n_1_230), .A1 (n_1_649), .A2 (n_1_647), .B1 (n_1_692), .B2 (n_1_618));
AOI221_X1 i_1_396 (.ZN (n_1_229), .A (n_1_230), .B1 (n_1_610), .B2 (n_1_487), .C1 (n_1_601), .C2 (n_1_505));
OAI211_X1 i_1_395 (.ZN (n_1_228), .A (n_1_231), .B (n_1_229), .C1 (n_1_707), .C2 (n_1_637));
OR4_X1 i_1_394 (.ZN (n_236), .A1 (n_1_234), .A2 (n_1_232), .A3 (n_1_242), .A4 (n_1_228));
OAI22_X1 i_1_393 (.ZN (n_1_227), .A1 (n_1_572), .A2 (n_1_247), .B1 (n_1_656), .B2 (n_1_584));
OAI22_X1 i_1_392 (.ZN (n_1_226), .A1 (n_1_713), .A2 (n_1_553), .B1 (n_1_647), .B2 (n_1_534));
NOR2_X2 i_1_391 (.ZN (n_1_225), .A1 (n_1_727), .A2 (n_1_722));
INV_X1 i_1_390 (.ZN (n_1_224), .A (n_1_225));
AOI22_X1 i_1_389 (.ZN (n_1_223), .A1 (n_1_564), .A2 (n_1_225), .B1 (n_1_702), .B2 (n_1_551));
OAI221_X1 i_1_388 (.ZN (n_1_222), .A (n_1_223), .B1 (n_1_707), .B2 (n_1_556), .C1 (n_1_724), .C2 (n_1_581));
OAI22_X1 i_1_387 (.ZN (n_1_221), .A1 (n_1_538), .A2 (n_1_486), .B1 (n_1_645), .B2 (n_1_547));
OAI22_X1 i_1_386 (.ZN (n_1_220), .A1 (n_1_704), .A2 (n_1_566), .B1 (n_1_692), .B2 (n_1_560));
AOI22_X1 i_1_385 (.ZN (n_1_219), .A1 (n_1_616), .A2 (n_1_532), .B1 (n_1_662), .B2 (n_1_542));
OAI221_X1 i_1_384 (.ZN (n_1_218), .A (n_1_219), .B1 (n_1_578), .B2 (n_1_516), .C1 (n_1_575), .C2 (n_1_504));
OR4_X1 i_1_383 (.ZN (n_1_217), .A1 (n_1_221), .A2 (n_1_220), .A3 (n_1_218), .A4 (n_1_222));
OR4_X1 i_1_382 (.ZN (n_235), .A1 (n_1_227), .A2 (n_1_226), .A3 (n_1_693), .A4 (n_1_217));
AOI22_X1 i_1_381 (.ZN (n_1_216), .A1 (drc_ipo_n19), .A2 (n_1_648), .B1 (n_1_662), .B2 (n_1_626));
OAI221_X1 i_1_380 (.ZN (n_1_215), .A (n_1_216), .B1 (n_1_701), .B2 (n_1_629), .C1 (n_1_600), .C2 (n_1_516));
OAI222_X1 i_1_379 (.ZN (n_1_214), .A1 (n_1_707), .A2 (n_1_605), .B1 (n_1_674), .B2 (n_1_617)
    , .C1 (n_1_649), .C2 (n_1_645));
AOI22_X1 i_1_378 (.ZN (n_1_213), .A1 (n_1_654), .A2 (n_1_225), .B1 (n_1_725), .B2 (n_1_685));
OAI221_X1 i_1_377 (.ZN (n_1_212), .A (n_1_213), .B1 (n_1_678), .B2 (n_1_504), .C1 (n_1_618), .C2 (n_1_247));
OAI22_X1 i_1_376 (.ZN (n_1_211), .A1 (n_1_596), .A2 (n_1_486), .B1 (n_1_713), .B2 (n_1_609));
OAI22_X1 i_1_375 (.ZN (n_1_210), .A1 (n_1_692), .A2 (n_1_637), .B1 (n_1_704), .B2 (n_1_670));
OR4_X1 i_1_374 (.ZN (n_1_209), .A1 (n_1_211), .A2 (n_1_210), .A3 (n_1_212), .A4 (n_1_214));
OR3_X1 i_1_373 (.ZN (n_234), .A1 (n_1_693), .A2 (n_1_215), .A3 (n_1_209));
OAI22_X1 i_1_372 (.ZN (n_1_208), .A1 (n_1_696), .A2 (n_1_563), .B1 (n_1_692), .B2 (n_1_556));
AOI221_X1 i_1_371 (.ZN (n_1_207), .A (n_1_208), .B1 (n_1_561), .B2 (n_1_248), .C1 (n_1_702), .C2 (n_1_582));
OAI211_X1 i_1_370 (.ZN (n_1_206), .A (n_1_698), .B (n_1_207), .C1 (n_1_617), .C2 (n_1_584));
OAI222_X1 i_1_369 (.ZN (n_1_205), .A1 (n_1_707), .A2 (n_1_553), .B1 (n_1_645), .B2 (n_1_534)
    , .C1 (n_1_704), .C2 (n_1_550));
AOI22_X1 i_1_368 (.ZN (n_1_204), .A1 (n_1_648), .A2 (n_1_579), .B1 (n_1_573), .B2 (n_1_225));
OAI221_X1 i_1_367 (.ZN (n_1_203), .A (n_1_204), .B1 (n_1_575), .B2 (n_1_516), .C1 (n_1_713), .C2 (n_1_538));
AOI22_X1 i_1_366 (.ZN (n_1_202), .A1 (n_1_725), .A2 (n_1_542), .B1 (n_1_662), .B2 (n_1_548));
OAI221_X1 i_1_365 (.ZN (n_1_201), .A (n_1_202), .B1 (n_1_566), .B2 (n_1_486), .C1 (n_1_531), .C2 (n_1_504));
OR4_X1 i_1_364 (.ZN (n_233), .A1 (n_1_203), .A2 (n_1_201), .A3 (n_1_205), .A4 (n_1_206));
AOI22_X1 i_1_363 (.ZN (n_1_200), .A1 (n_1_671), .A2 (n_1_487), .B1 (n_1_702), .B2 (n_1_685));
OAI221_X1 i_1_362 (.ZN (n_1_199), .A (n_1_200), .B1 (n_1_678), .B2 (n_1_516), .C1 (n_1_674), .C2 (n_1_504));
AOI21_X1 i_1_361 (.ZN (n_1_198), .A (n_1_699), .B1 (n_1_662), .B2 (n_1_650));
OAI221_X1 i_1_360 (.ZN (n_1_197), .A (n_1_198), .B1 (n_1_618), .B2 (n_1_224), .C1 (n_1_696), .C2 (n_1_653));
AOI22_X1 i_1_359 (.ZN (n_1_196), .A1 (n_1_712), .A2 (n_1_597), .B1 (n_1_708), .B2 (n_1_610));
OAI221_X1 i_1_358 (.ZN (n_1_195), .A (n_1_196), .B1 (n_1_692), .B2 (n_1_605), .C1 (n_1_704), .C2 (n_1_629));
AOI22_X1 i_1_357 (.ZN (n_1_194), .A1 (drc_ipo_n19), .A2 (n_1_646), .B1 (n_1_638), .B2 (n_1_248));
OAI221_X1 i_1_356 (.ZN (n_1_193), .A (n_1_194), .B1 (n_1_647), .B2 (n_1_600), .C1 (n_1_724), .C2 (n_1_625));
OR4_X1 i_1_355 (.ZN (n_232), .A1 (n_1_199), .A2 (n_1_197), .A3 (n_1_195), .A4 (n_1_193));
AOI22_X1 i_1_354 (.ZN (n_1_192), .A1 (n_1_708), .A2 (n_1_539), .B1 (n_1_648), .B2 (n_1_576));
OAI221_X1 i_1_353 (.ZN (n_1_191), .A (n_1_192), .B1 (n_1_531), .B2 (n_1_516), .C1 (n_1_701), .C2 (n_1_541));
AOI22_X1 i_1_352 (.ZN (n_1_190), .A1 (n_1_561), .A2 (n_1_225), .B1 (n_1_712), .B2 (n_1_567));
OAI221_X1 i_1_351 (.ZN (n_1_189), .A (n_1_190), .B1 (n_1_645), .B2 (n_1_578), .C1 (n_1_584), .C2 (n_1_504));
OAI22_X1 i_1_350 (.ZN (n_1_188), .A1 (n_1_692), .A2 (n_1_553), .B1 (n_1_704), .B2 (n_1_581));
INV_X1 i_1_349 (.ZN (n_1_187), .A (n_1_188));
OAI221_X1 i_1_348 (.ZN (n_1_186), .A (n_1_187), .B1 (n_1_550), .B2 (n_1_486), .C1 (hfn_ipo_n15), .C2 (n_1_563));
AOI22_X1 i_1_347 (.ZN (n_1_185), .A1 (n_1_557), .A2 (n_1_248), .B1 (n_1_725), .B2 (n_1_548));
OAI221_X1 i_1_346 (.ZN (n_1_184), .A (n_1_185), .B1 (n_1_696), .B2 (n_1_572), .C1 (n_1_661), .C2 (n_1_534));
OR4_X1 i_1_345 (.ZN (n_231), .A1 (n_1_191), .A2 (n_1_189), .A3 (n_1_186), .A4 (n_1_184));
AOI22_X1 i_1_344 (.ZN (n_1_183), .A1 (n_1_675), .A2 (n_1_517), .B1 (drc_ipo_n19), .B2 (n_1_662));
OAI221_X1 i_1_343 (.ZN (n_1_182), .A (n_1_183), .B1 (n_1_645), .B2 (n_1_600), .C1 (n_1_692), .C2 (n_1_609));
AOI22_X1 i_1_342 (.ZN (n_1_181), .A1 (n_1_606), .A2 (n_1_248), .B1 (n_1_638), .B2 (n_1_225));
OAI221_X1 i_1_341 (.ZN (n_1_180), .A (n_1_181), .B1 (n_1_707), .B2 (n_1_596), .C1 (n_1_701), .C2 (n_1_625));
OAI222_X1 i_1_340 (.ZN (n_1_179), .A1 (n_1_713), .A2 (n_1_670), .B1 (n_1_704), .B2 (n_1_684)
    , .C1 (hfn_ipo_n15), .C2 (n_1_653));
AOI22_X1 i_1_339 (.ZN (n_1_178), .A1 (n_1_679), .A2 (n_1_648), .B1 (n_1_630), .B2 (n_1_487));
OAI221_X1 i_1_338 (.ZN (n_1_177), .A (n_1_178), .B1 (n_1_696), .B2 (n_1_618), .C1 (n_1_724), .C2 (n_1_649));
OR4_X1 i_1_337 (.ZN (n_230), .A1 (n_1_182), .A2 (n_1_180), .A3 (n_1_179), .A4 (n_1_177));
OAI22_X1 i_1_336 (.ZN (n_1_176), .A1 (n_1_724), .A2 (n_1_534), .B1 (n_1_692), .B2 (n_1_538));
INV_X1 i_1_335 (.ZN (n_1_175), .A (n_1_176));
OAI221_X1 i_1_334 (.ZN (n_1_174), .A (n_1_175), .B1 (n_1_701), .B2 (n_1_547), .C1 (n_1_661), .C2 (n_1_578));
AOI22_X1 i_1_333 (.ZN (n_1_173), .A1 (n_1_708), .A2 (n_1_567), .B1 (n_1_582), .B2 (n_1_487));
OAI221_X1 i_1_332 (.ZN (n_1_172), .A (n_1_173), .B1 (n_1_713), .B2 (n_1_550), .C1 (n_1_584), .C2 (n_1_516));
OAI222_X1 i_1_331 (.ZN (n_1_171), .A1 (n_1_556), .A2 (n_1_224), .B1 (n_1_553), .B2 (n_1_247)
    , .C1 (n_1_704), .C2 (n_1_541));
AOI22_X1 i_1_330 (.ZN (n_1_170), .A1 (hfn_ipo_n14), .A2 (n_1_573), .B1 (n_1_648), .B2 (n_1_532));
OAI221_X1 i_1_329 (.ZN (n_1_169), .A (n_1_170), .B1 (n_1_645), .B2 (n_1_575), .C1 (n_1_696), .C2 (n_1_560));
OR4_X1 i_1_328 (.ZN (n_229), .A1 (n_1_174), .A2 (n_1_172), .A3 (n_1_171), .A4 (n_1_169));
OAI22_X1 i_1_327 (.ZN (n_1_168), .A1 (n_1_724), .A2 (n_1_664), .B1 (n_1_713), .B2 (n_1_629));
AOI221_X1 i_1_326 (.ZN (n_1_167), .A (n_1_168), .B1 (hfn_ipo_n13), .B2 (n_1_619), .C1 (n_1_697), .C2 (n_1_638));
OAI221_X1 i_1_325 (.ZN (n_1_166), .A (n_1_167), .B1 (n_1_704), .B2 (n_1_625), .C1 (n_1_701), .C2 (n_1_649));
AOI22_X1 i_1_324 (.ZN (n_1_165), .A1 (n_1_662), .A2 (n_1_601), .B1 (n_1_675), .B2 (n_1_648));
OAI221_X1 i_1_323 (.ZN (n_1_164), .A (n_1_165), .B1 (n_1_692), .B2 (n_1_596), .C1 (n_1_707), .C2 (n_1_670));
OAI22_X1 i_1_322 (.ZN (n_1_163), .A1 (n_1_684), .A2 (n_1_486), .B1 (n_1_609), .B2 (n_1_247));
OAI22_X1 i_1_321 (.ZN (n_1_162), .A1 (n_1_605), .A2 (n_1_224), .B1 (n_1_678), .B2 (n_1_645));
OR4_X1 i_1_320 (.ZN (n_228), .A1 (n_1_163), .A2 (n_1_162), .A3 (n_1_164), .A4 (n_1_166));
OAI22_X1 i_1_319 (.ZN (n_1_161), .A1 (n_1_696), .A2 (n_1_556), .B1 (n_1_707), .B2 (n_1_550));
AOI221_X1 i_1_318 (.ZN (n_1_160), .A (n_1_161), .B1 (n_1_554), .B2 (n_1_225), .C1 (n_1_712), .C2 (n_1_582));
OAI221_X1 i_1_317 (.ZN (n_1_159), .A (n_1_160), .B1 (n_1_701), .B2 (n_1_534), .C1 (n_1_647), .C2 (n_1_584));
AOI22_X1 i_1_316 (.ZN (n_1_158), .A1 (n_1_542), .A2 (n_1_487), .B1 (n_1_662), .B2 (n_1_576));
OAI221_X1 i_1_315 (.ZN (n_1_157), .A (n_1_158), .B1 (n_1_692), .B2 (n_1_566), .C1 (hfn_ipo_n15), .C2 (n_1_560));
OAI22_X1 i_1_314 (.ZN (n_1_156), .A1 (n_1_724), .A2 (n_1_578), .B1 (n_1_704), .B2 (n_1_547));
OAI22_X1 i_1_313 (.ZN (n_1_155), .A1 (n_1_538), .A2 (n_1_247), .B1 (n_1_645), .B2 (n_1_531));
OR4_X1 i_1_312 (.ZN (n_227), .A1 (n_1_156), .A2 (n_1_155), .A3 (n_1_157), .A4 (n_1_159));
OAI22_X1 i_1_311 (.ZN (n_1_154), .A1 (n_1_674), .A2 (n_1_645), .B1 (n_1_692), .B2 (n_1_670));
AOI221_X1 i_1_310 (.ZN (n_1_153), .A (n_1_154), .B1 (n_1_626), .B2 (n_1_487), .C1 (n_1_725), .C2 (n_1_601));
OAI221_X1 i_1_309 (.ZN (n_1_152), .A (n_1_153), .B1 (hfn_ipo_n15), .B2 (n_1_637), .C1 (n_1_696), .C2 (n_1_605));
OAI222_X1 i_1_308 (.ZN (n_1_151), .A1 (n_1_704), .A2 (n_1_649), .B1 (n_1_701), .B2 (n_1_664)
    , .C1 (n_1_678), .C2 (n_1_661));
OAI22_X1 i_1_307 (.ZN (n_1_150), .A1 (n_1_596), .A2 (n_1_247), .B1 (n_1_707), .B2 (n_1_629));
OAI22_X1 i_1_306 (.ZN (n_1_149), .A1 (n_1_713), .A2 (n_1_684), .B1 (n_1_609), .B2 (n_1_224));
OR4_X1 i_1_305 (.ZN (n_226), .A1 (n_1_150), .A2 (n_1_149), .A3 (n_1_151), .A4 (n_1_152));
OAI22_X1 i_1_304 (.ZN (n_1_148), .A1 (n_1_547), .A2 (n_1_486), .B1 (n_1_696), .B2 (n_1_553));
AOI221_X1 i_1_303 (.ZN (n_1_147), .A (n_1_148), .B1 (n_1_567), .B2 (n_1_248), .C1 (n_1_662), .C2 (n_1_532));
OAI221_X1 i_1_302 (.ZN (n_1_146), .A (n_1_147), .B1 (n_1_704), .B2 (n_1_534), .C1 (n_1_645), .C2 (n_1_584));
OAI222_X1 i_1_301 (.ZN (n_1_145), .A1 (n_1_701), .A2 (n_1_578), .B1 (n_1_724), .B2 (n_1_575)
    , .C1 (n_1_713), .C2 (n_1_541));
AOI22_X1 i_1_300 (.ZN (n_1_144), .A1 (n_1_708), .A2 (n_1_582), .B1 (hfn_ipo_n13), .B2 (n_1_557));
OAI221_X1 i_1_299 (.ZN (n_1_143), .A (n_1_144), .B1 (n_1_692), .B2 (n_1_550), .C1 (n_1_538), .C2 (n_1_224));
OR3_X1 i_1_298 (.ZN (n_225), .A1 (n_1_145), .A2 (n_1_143), .A3 (n_1_146));
AOI22_X1 i_1_297 (.ZN (n_1_142), .A1 (n_1_697), .A2 (n_1_610), .B1 (n_1_725), .B2 (n_1_679));
OAI221_X1 i_1_296 (.ZN (n_1_141), .A (n_1_142), .B1 (n_1_649), .B2 (n_1_486), .C1 (n_1_713), .C2 (n_1_625));
OAI22_X1 i_1_295 (.ZN (n_1_140), .A1 (n_1_701), .A2 (n_1_600), .B1 (n_1_704), .B2 (n_1_664));
INV_X1 i_1_294 (.ZN (n_1_139), .A (n_1_140));
OAI221_X1 i_1_293 (.ZN (n_1_138), .A (n_1_139), .B1 (n_1_670), .B2 (n_1_247), .C1 (hfn_ipo_n15), .C2 (n_1_605));
OAI22_X1 i_1_292 (.ZN (n_1_137), .A1 (n_1_692), .A2 (n_1_629), .B1 (n_1_674), .B2 (n_1_661));
OAI22_X1 i_1_291 (.ZN (n_1_136), .A1 (n_1_596), .A2 (n_1_224), .B1 (n_1_707), .B2 (n_1_684));
OR4_X1 i_1_290 (.ZN (n_224), .A1 (n_1_137), .A2 (n_1_136), .A3 (n_1_138), .A4 (n_1_141));
AOI22_X1 i_1_289 (.ZN (n_1_135), .A1 (n_1_567), .A2 (n_1_225), .B1 (n_1_697), .B2 (n_1_539));
OAI221_X1 i_1_288 (.ZN (n_1_134), .A (n_1_135), .B1 (n_1_534), .B2 (n_1_486), .C1 (n_1_701), .C2 (n_1_575));
OAI22_X1 i_1_287 (.ZN (n_1_133), .A1 (n_1_707), .A2 (n_1_541), .B1 (n_1_692), .B2 (n_1_581));
INV_X1 i_1_286 (.ZN (n_1_132), .A (n_1_133));
OAI221_X1 i_1_285 (.ZN (n_1_131), .A (n_1_132), .B1 (n_1_704), .B2 (n_1_578), .C1 (hfn_ipo_n16), .C2 (n_1_553));
OAI22_X1 i_1_284 (.ZN (n_1_130), .A1 (n_1_724), .A2 (n_1_531), .B1 (n_1_661), .B2 (n_1_584));
OAI22_X1 i_1_283 (.ZN (n_1_129), .A1 (n_1_550), .A2 (n_1_247), .B1 (n_1_713), .B2 (n_1_547));
OR4_X1 i_1_282 (.ZN (n_223), .A1 (n_1_130), .A2 (n_1_129), .A3 (n_1_131), .A4 (n_1_134));
OAI222_X1 i_1_281 (.ZN (n_1_128), .A1 (n_1_704), .A2 (n_1_600), .B1 (n_1_670), .B2 (n_1_224)
    , .C1 (n_1_696), .C2 (n_1_596));
OAI22_X1 i_1_280 (.ZN (n_1_127), .A1 (n_1_629), .A2 (n_1_247), .B1 (n_1_692), .B2 (n_1_684));
INV_X1 i_1_279 (.ZN (n_1_126), .A (n_1_127));
OAI221_X1 i_1_278 (.ZN (n_1_125), .A (n_1_126), .B1 (n_1_701), .B2 (n_1_678), .C1 (n_1_707), .C2 (n_1_625));
OAI22_X1 i_1_277 (.ZN (n_1_124), .A1 (hfn_ipo_n16), .A2 (n_1_609), .B1 (n_1_664), .B2 (n_1_486));
OAI22_X1 i_1_276 (.ZN (n_1_123), .A1 (n_1_724), .A2 (n_1_674), .B1 (n_1_713), .B2 (n_1_649));
OR4_X1 i_1_275 (.ZN (n_222), .A1 (n_1_124), .A2 (n_1_123), .A3 (n_1_125), .A4 (n_1_128));
OAI222_X1 i_1_274 (.ZN (n_1_122), .A1 (n_1_704), .A2 (n_1_575), .B1 (n_1_692), .B2 (n_1_541)
    , .C1 (n_1_701), .C2 (n_1_531));
AOI22_X1 i_1_273 (.ZN (n_1_121), .A1 (n_1_708), .A2 (n_1_548), .B1 (n_1_579), .B2 (n_1_487));
OAI221_X1 i_1_272 (.ZN (n_1_120), .A (n_1_121), .B1 (n_1_713), .B2 (n_1_534), .C1 (hfn_ipo_n15), .C2 (n_1_538));
OAI22_X1 i_1_271 (.ZN (n_1_119), .A1 (n_1_696), .A2 (n_1_566), .B1 (n_1_724), .B2 (n_1_584));
OAI22_X1 i_1_270 (.ZN (n_1_118), .A1 (n_1_550), .A2 (n_1_224), .B1 (n_1_581), .B2 (n_1_247));
OR4_X1 i_1_269 (.ZN (n_221), .A1 (n_1_119), .A2 (n_1_118), .A3 (n_1_120), .A4 (n_1_122));
OAI22_X1 i_1_268 (.ZN (n_1_117), .A1 (n_1_684), .A2 (n_1_247), .B1 (n_1_600), .B2 (n_1_486));
OAI22_X1 i_1_267 (.ZN (n_1_116), .A1 (n_1_629), .A2 (n_1_224), .B1 (n_1_704), .B2 (n_1_678));
OAI22_X1 i_1_266 (.ZN (n_1_115), .A1 (n_1_692), .A2 (n_1_625), .B1 (n_1_701), .B2 (n_1_674));
AOI221_X1 i_1_265 (.ZN (n_1_114), .A (n_1_115), .B1 (n_1_712), .B2 (drc_ipo_n19), .C1 (n_1_708), .C2 (n_1_650));
OAI221_X1 i_1_264 (.ZN (n_1_113), .A (n_1_114), .B1 (hfn_ipo_n15), .B2 (n_1_596), .C1 (n_1_696), .C2 (n_1_670));
OR3_X1 i_1_263 (.ZN (n_220), .A1 (n_1_117), .A2 (n_1_116), .A3 (n_1_113));
OAI22_X1 i_1_262 (.ZN (n_1_112), .A1 (n_1_575), .A2 (n_1_486), .B1 (n_1_704), .B2 (n_1_531));
OAI22_X1 i_1_261 (.ZN (n_1_111), .A1 (n_1_713), .A2 (n_1_578), .B1 (hfn_ipo_n15), .B2 (n_1_566));
OAI22_X1 i_1_260 (.ZN (n_1_110), .A1 (n_1_581), .A2 (n_1_224), .B1 (n_1_692), .B2 (n_1_547));
AOI221_X1 i_1_259 (.ZN (n_1_109), .A (n_1_110), .B1 (n_1_708), .B2 (n_1_535), .C1 (n_1_542), .C2 (n_1_248));
OAI221_X1 i_1_258 (.ZN (n_1_108), .A (n_1_109), .B1 (n_1_701), .B2 (n_1_584), .C1 (n_1_696), .C2 (n_1_550));
OR3_X1 i_1_257 (.ZN (n_219), .A1 (n_1_112), .A2 (n_1_111), .A3 (n_1_108));
OAI22_X1 i_1_256 (.ZN (n_1_107), .A1 (hfn_ipo_n15), .A2 (n_1_670), .B1 (n_1_692), .B2 (n_1_649));
OAI22_X1 i_1_255 (.ZN (n_1_106), .A1 (n_1_704), .A2 (n_1_674), .B1 (n_1_696), .B2 (n_1_629));
AOI221_X1 i_1_254 (.ZN (n_1_105), .A (n_1_106), .B1 (n_1_626), .B2 (n_1_248), .C1 (n_1_679), .C2 (n_1_487));
OAI221_X1 i_1_253 (.ZN (n_1_104), .A (n_1_105), .B1 (n_1_684), .B2 (n_1_224), .C1 (n_1_713), .C2 (n_1_600));
AOI211_X1 i_1_252 (.ZN (n_1_103), .A (n_1_107), .B (n_1_104), .C1 (n_1_708), .C2 (drc_ipo_n19));
INV_X1 i_1_251 (.ZN (n_218), .A (n_1_103));
OAI22_X1 i_1_250 (.ZN (n_1_102), .A1 (n_1_692), .A2 (n_1_534), .B1 (n_1_707), .B2 (n_1_578));
OAI22_X1 i_1_249 (.ZN (n_1_101), .A1 (n_1_696), .A2 (n_1_581), .B1 (n_1_547), .B2 (n_1_247));
AOI221_X1 i_1_248 (.ZN (n_1_100), .A (n_1_101), .B1 (n_1_712), .B2 (n_1_576), .C1 (hfn_ipo_n13), .C2 (n_1_551));
OAI221_X1 i_1_247 (.ZN (n_1_99), .A (n_1_100), .B1 (n_1_531), .B2 (n_1_486), .C1 (n_1_704), .C2 (n_1_584));
AOI211_X1 i_1_246 (.ZN (n_1_98), .A (n_1_102), .B (n_1_99), .C1 (n_1_542), .C2 (n_1_225));
INV_X1 i_1_245 (.ZN (n_217), .A (n_1_98));
OAI22_X1 i_1_244 (.ZN (n_1_97), .A1 (n_1_649), .A2 (n_1_247), .B1 (n_1_625), .B2 (n_1_224));
OAI22_X1 i_1_243 (.ZN (n_1_96), .A1 (hfn_ipo_n16), .A2 (n_1_629), .B1 (n_1_696), .B2 (n_1_684));
AOI22_X1 i_1_242 (.ZN (n_1_95), .A1 (n_1_675), .A2 (n_1_487), .B1 (n_1_712), .B2 (n_1_679));
OAI221_X1 i_1_241 (.ZN (n_1_94), .A (n_1_95), .B1 (n_1_692), .B2 (n_1_664), .C1 (n_1_707), .C2 (n_1_600));
OR3_X1 i_1_240 (.ZN (n_216), .A1 (n_1_97), .A2 (n_1_96), .A3 (n_1_94));
OAI22_X1 i_1_239 (.ZN (n_1_93), .A1 (n_1_547), .A2 (n_1_224), .B1 (n_1_696), .B2 (n_1_541));
OAI22_X1 i_1_238 (.ZN (n_1_92), .A1 (n_1_534), .A2 (n_1_247), .B1 (n_1_692), .B2 (n_1_578));
AOI22_X1 i_1_237 (.ZN (n_1_91), .A1 (hfn_ipo_n13), .A2 (n_1_582), .B1 (n_1_708), .B2 (n_1_576));
OAI221_X1 i_1_236 (.ZN (n_1_90), .A (n_1_91), .B1 (n_1_713), .B2 (n_1_531), .C1 (n_1_584), .C2 (n_1_486));
OR3_X1 i_1_235 (.ZN (n_215), .A1 (n_1_93), .A2 (n_1_92), .A3 (n_1_90));
AOI22_X1 i_1_234 (.ZN (n_1_89), .A1 (n_1_712), .A2 (n_1_675), .B1 (hfn_ipo_n13), .B2 (n_1_685));
OAI22_X1 i_1_233 (.ZN (n_1_88), .A1 (n_1_692), .A2 (n_1_600), .B1 (n_1_664), .B2 (n_1_247));
AOI221_X1 i_1_232 (.ZN (n_1_87), .A (n_1_88), .B1 (n_1_650), .B2 (n_1_225), .C1 (n_1_708), .C2 (n_1_679));
OAI211_X1 i_1_231 (.ZN (n_214), .A (n_1_89), .B (n_1_87), .C1 (n_1_696), .C2 (n_1_625));
OAI22_X1 i_1_230 (.ZN (n_1_86), .A1 (n_1_692), .A2 (n_1_575), .B1 (n_1_707), .B2 (n_1_531));
INV_X1 i_1_229 (.ZN (n_1_85), .A (n_1_86));
OAI22_X1 i_1_228 (.ZN (n_1_84), .A1 (hfn_ipo_n15), .A2 (n_1_541), .B1 (n_1_713), .B2 (n_1_584));
AOI221_X1 i_1_227 (.ZN (n_1_83), .A (n_1_84), .B1 (n_1_697), .B2 (n_1_548), .C1 (n_1_579), .C2 (n_1_248));
OAI211_X1 i_1_226 (.ZN (n_213), .A (n_1_85), .B (n_1_83), .C1 (n_1_534), .C2 (n_1_224));
OAI22_X1 i_1_225 (.ZN (n_1_82), .A1 (n_1_692), .A2 (n_1_678), .B1 (hfn_ipo_n15), .B2 (n_1_625));
AOI221_X1 i_1_224 (.ZN (n_1_81), .A (n_1_82), .B1 (drc_ipo_n19), .B2 (n_1_225), .C1 (n_1_697), .C2 (n_1_650));
OAI221_X1 i_1_223 (.ZN (n_212), .A (n_1_81), .B1 (n_1_707), .B2 (n_1_674), .C1 (n_1_600), .C2 (n_1_247));
OAI22_X1 i_1_222 (.ZN (n_1_80), .A1 (n_1_692), .A2 (n_1_531), .B1 (n_1_578), .B2 (n_1_224));
AOI221_X1 i_1_221 (.ZN (n_1_79), .A (n_1_80), .B1 (n_1_576), .B2 (n_1_248), .C1 (n_1_697), .C2 (n_1_535));
OAI221_X1 i_1_220 (.ZN (n_211), .A (n_1_79), .B1 (hfn_ipo_n15), .B2 (n_1_547), .C1 (n_1_707), .C2 (n_1_584));
OAI22_X1 i_1_219 (.ZN (n_1_78), .A1 (n_1_692), .A2 (n_1_674), .B1 (n_1_678), .B2 (n_1_247));
AOI21_X1 i_1_218 (.ZN (n_1_77), .A (n_1_78), .B1 (n_1_697), .B2 (drc_ipo_n19));
OAI221_X1 i_1_217 (.ZN (n_210), .A (n_1_77), .B1 (n_1_600), .B2 (n_1_224), .C1 (hfn_ipo_n15), .C2 (n_1_649));
AOI222_X1 i_1_216 (.ZN (n_1_76), .A1 (hfn_ipo_n13), .A2 (n_1_535), .B1 (n_1_697), .B2 (n_1_579)
    , .C1 (n_1_532), .C2 (n_1_248));
OAI221_X1 i_1_215 (.ZN (n_209), .A (n_1_76), .B1 (n_1_575), .B2 (n_1_224), .C1 (n_1_692), .C2 (n_1_584));
AOI22_X1 i_1_214 (.ZN (n_1_75), .A1 (hfn_ipo_n13), .A2 (drc_ipo_n19), .B1 (n_1_697), .B2 (n_1_601));
OAI221_X1 i_1_213 (.ZN (n_208), .A (n_1_75), .B1 (n_1_674), .B2 (n_1_247), .C1 (n_1_678), .C2 (n_1_224));
AOI22_X1 i_1_212 (.ZN (n_1_74), .A1 (n_1_697), .A2 (n_1_576), .B1 (n_1_532), .B2 (n_1_225));
OAI221_X1 i_1_211 (.ZN (n_207), .A (n_1_74), .B1 (hfn_ipo_n15), .B2 (n_1_578), .C1 (n_1_584), .C2 (n_1_247));
OAI222_X1 i_1_210 (.ZN (n_206), .A1 (n_1_674), .A2 (n_1_224), .B1 (n_1_696), .B2 (n_1_678)
    , .C1 (hfn_ipo_n16), .C2 (n_1_600));
OAI222_X1 i_1_209 (.ZN (n_205), .A1 (n_1_696), .A2 (n_1_531), .B1 (n_1_584), .B2 (n_1_224)
    , .C1 (hfn_ipo_n16), .C2 (n_1_575));
OAI22_X1 i_1_208 (.ZN (n_204), .A1 (n_1_696), .A2 (n_1_674), .B1 (hfn_ipo_n16), .B2 (n_1_678));
OAI22_X1 i_1_207 (.ZN (n_203), .A1 (n_1_696), .A2 (n_1_584), .B1 (hfn_ipo_n15), .B2 (n_1_531));
NOR2_X1 i_1_206 (.ZN (n_202), .A1 (hfn_ipo_n15), .A2 (n_1_674));
NOR2_X1 i_1_205 (.ZN (n_201), .A1 (hfn_ipo_n15), .A2 (n_1_584));
NAND2_X2 i_1_204 (.ZN (n_1_73), .A1 (n_1_924), .A2 (b[0]));
NAND2_X2 i_1_203 (.ZN (n_1_72), .A1 (b[1]), .A2 (n_1_923));
NAND2_X2 i_1_202 (.ZN (n_1_71), .A1 (b[1]), .A2 (b[0]));
OAI222_X1 i_1_201 (.ZN (n_1_70), .A1 (n_1_920), .A2 (n_1_72), .B1 (n_1_921), .B2 (n_1_71)
    , .C1 (n_1_890), .C2 (n_1_73));
NAND2_X4 i_1_200 (.ZN (n_1_69), .A1 (hfn_ipo_n13), .A2 (n_1_70));
OAI21_X1 i_1_199 (.ZN (n_200), .A (n_1_69), .B1 (n_1_858), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_198 (.ZN (n_199), .A (n_1_69), .B1 (n_1_857), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_197 (.ZN (n_198), .A (n_1_69), .B1 (n_1_856), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_196 (.ZN (n_197), .A (n_1_69), .B1 (n_1_855), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_195 (.ZN (n_196), .A (n_1_69), .B1 (n_1_854), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_194 (.ZN (n_195), .A (n_1_69), .B1 (n_1_853), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_193 (.ZN (n_194), .A (n_1_69), .B1 (n_1_852), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_192 (.ZN (n_193), .A (n_1_69), .B1 (n_1_851), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_191 (.ZN (n_192), .A (n_1_69), .B1 (n_1_850), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_190 (.ZN (n_191), .A (n_1_69), .B1 (n_1_849), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_189 (.ZN (n_190), .A (n_1_69), .B1 (n_1_848), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_188 (.ZN (n_189), .A (n_1_69), .B1 (n_1_847), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_187 (.ZN (n_188), .A (n_1_69), .B1 (n_1_846), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_186 (.ZN (n_187), .A (n_1_69), .B1 (n_1_845), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_185 (.ZN (n_186), .A (n_1_69), .B1 (n_1_844), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_184 (.ZN (n_185), .A (n_1_69), .B1 (n_1_843), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_183 (.ZN (n_184), .A (n_1_69), .B1 (n_1_842), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_182 (.ZN (n_183), .A (n_1_69), .B1 (n_1_841), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_181 (.ZN (n_182), .A (n_1_69), .B1 (n_1_840), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_180 (.ZN (n_181), .A (n_1_69), .B1 (n_1_839), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_179 (.ZN (n_180), .A (n_1_69), .B1 (n_1_838), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_178 (.ZN (n_179), .A (n_1_69), .B1 (n_1_837), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_177 (.ZN (n_178), .A (n_1_69), .B1 (n_1_836), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_176 (.ZN (n_177), .A (n_1_69), .B1 (n_1_835), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_175 (.ZN (n_176), .A (n_1_69), .B1 (n_1_834), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_174 (.ZN (n_175), .A (n_1_69), .B1 (n_1_833), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_173 (.ZN (n_174), .A (n_1_69), .B1 (n_1_832), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_172 (.ZN (n_173), .A (n_1_69), .B1 (n_1_831), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_171 (.ZN (n_172), .A (n_1_69), .B1 (n_1_830), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_170 (.ZN (n_171), .A (n_1_69), .B1 (n_1_829), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_169 (.ZN (n_170), .A (n_1_69), .B1 (n_1_828), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_168 (.ZN (n_169), .A (n_1_69), .B1 (n_1_827), .B2 (hfn_ipo_n14));
OAI21_X1 i_1_167 (.ZN (n_168), .A (n_1_69), .B1 (n_1_826), .B2 (hfn_ipo_n14));
OAI222_X1 i_1_166 (.ZN (n_1_68), .A1 (n_1_889), .A2 (n_1_73), .B1 (n_1_919), .B2 (n_1_72)
    , .C1 (n_1_920), .C2 (n_1_71));
INV_X1 i_1_165 (.ZN (n_1_67), .A (n_1_68));
OAI22_X1 i_1_164 (.ZN (n_167), .A1 (n_1_825), .A2 (hfn_ipo_n14), .B1 (hfn_ipo_n16), .B2 (n_1_67));
OAI222_X1 i_1_163 (.ZN (n_1_66), .A1 (n_1_888), .A2 (n_1_73), .B1 (n_1_918), .B2 (n_1_72)
    , .C1 (n_1_919), .C2 (n_1_71));
INV_X1 i_1_162 (.ZN (n_1_65), .A (n_1_66));
OAI22_X1 i_1_161 (.ZN (n_166), .A1 (n_1_824), .A2 (hfn_ipo_n14), .B1 (hfn_ipo_n16), .B2 (n_1_65));
OAI222_X1 i_1_160 (.ZN (n_1_64), .A1 (n_1_887), .A2 (n_1_73), .B1 (n_1_917), .B2 (n_1_72)
    , .C1 (n_1_918), .C2 (n_1_71));
INV_X1 i_1_159 (.ZN (n_1_63), .A (n_1_64));
OAI22_X1 i_1_158 (.ZN (n_165), .A1 (n_1_823), .A2 (hfn_ipo_n14), .B1 (hfn_ipo_n16), .B2 (n_1_63));
OAI222_X1 i_1_157 (.ZN (n_1_62), .A1 (n_1_886), .A2 (n_1_73), .B1 (n_1_916), .B2 (n_1_72)
    , .C1 (n_1_917), .C2 (n_1_71));
INV_X1 i_1_156 (.ZN (n_1_61), .A (n_1_62));
OAI22_X1 i_1_155 (.ZN (n_164), .A1 (n_1_822), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_61));
OAI222_X1 i_1_154 (.ZN (n_1_60), .A1 (n_1_885), .A2 (n_1_73), .B1 (n_1_915), .B2 (n_1_72)
    , .C1 (n_1_916), .C2 (n_1_71));
INV_X1 i_1_153 (.ZN (n_1_59), .A (n_1_60));
OAI22_X1 i_1_152 (.ZN (n_163), .A1 (n_1_821), .A2 (hfn_ipo_n14), .B1 (hfn_ipo_n16), .B2 (n_1_59));
OAI222_X1 i_1_151 (.ZN (n_1_58), .A1 (n_1_884), .A2 (n_1_73), .B1 (n_1_914), .B2 (n_1_72)
    , .C1 (n_1_915), .C2 (n_1_71));
INV_X1 i_1_150 (.ZN (n_1_57), .A (n_1_58));
OAI22_X1 i_1_149 (.ZN (n_162), .A1 (n_1_820), .A2 (hfn_ipo_n14), .B1 (hfn_ipo_n16), .B2 (n_1_57));
OAI222_X1 i_1_148 (.ZN (n_1_56), .A1 (n_1_883), .A2 (n_1_73), .B1 (n_1_913), .B2 (n_1_72)
    , .C1 (n_1_914), .C2 (n_1_71));
INV_X1 i_1_147 (.ZN (n_1_55), .A (n_1_56));
OAI22_X1 i_1_146 (.ZN (n_161), .A1 (n_1_819), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_55));
OAI222_X1 i_1_145 (.ZN (n_1_54), .A1 (n_1_882), .A2 (n_1_73), .B1 (n_1_912), .B2 (n_1_72)
    , .C1 (n_1_913), .C2 (n_1_71));
INV_X1 i_1_144 (.ZN (n_1_53), .A (n_1_54));
OAI22_X1 i_1_143 (.ZN (n_160), .A1 (n_1_818), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_53));
OAI222_X1 i_1_142 (.ZN (n_1_52), .A1 (n_1_881), .A2 (n_1_73), .B1 (n_1_911), .B2 (n_1_72)
    , .C1 (n_1_912), .C2 (n_1_71));
INV_X1 i_1_141 (.ZN (n_1_51), .A (n_1_52));
OAI22_X1 i_1_140 (.ZN (n_159), .A1 (n_1_817), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_51));
OAI222_X1 i_1_139 (.ZN (n_1_50), .A1 (n_1_880), .A2 (n_1_73), .B1 (n_1_910), .B2 (n_1_72)
    , .C1 (n_1_911), .C2 (n_1_71));
INV_X1 i_1_138 (.ZN (n_1_49), .A (n_1_50));
OAI22_X1 i_1_137 (.ZN (n_158), .A1 (n_1_816), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_49));
OAI222_X1 i_1_136 (.ZN (n_1_48), .A1 (n_1_879), .A2 (n_1_73), .B1 (n_1_909), .B2 (n_1_72)
    , .C1 (n_1_910), .C2 (n_1_71));
INV_X1 i_1_135 (.ZN (n_1_47), .A (n_1_48));
OAI22_X1 i_1_134 (.ZN (n_157), .A1 (n_1_815), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_47));
OAI222_X1 i_1_133 (.ZN (n_1_46), .A1 (n_1_878), .A2 (n_1_73), .B1 (n_1_908), .B2 (n_1_72)
    , .C1 (n_1_909), .C2 (n_1_71));
INV_X1 i_1_132 (.ZN (n_1_45), .A (n_1_46));
OAI22_X1 i_1_131 (.ZN (n_156), .A1 (n_1_814), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_45));
OAI222_X1 i_1_130 (.ZN (n_1_44), .A1 (n_1_877), .A2 (n_1_73), .B1 (n_1_907), .B2 (n_1_72)
    , .C1 (n_1_908), .C2 (n_1_71));
INV_X1 i_1_129 (.ZN (n_1_43), .A (n_1_44));
OAI22_X1 i_1_128 (.ZN (n_155), .A1 (n_1_813), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_43));
OAI222_X1 i_1_127 (.ZN (n_1_42), .A1 (n_1_876), .A2 (n_1_73), .B1 (n_1_906), .B2 (n_1_72)
    , .C1 (n_1_907), .C2 (n_1_71));
INV_X1 i_1_126 (.ZN (n_1_41), .A (n_1_42));
OAI22_X1 i_1_125 (.ZN (n_154), .A1 (n_1_812), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_41));
OAI222_X1 i_1_124 (.ZN (n_1_40), .A1 (n_1_875), .A2 (n_1_73), .B1 (n_1_905), .B2 (n_1_72)
    , .C1 (n_1_906), .C2 (n_1_71));
INV_X1 i_1_123 (.ZN (n_1_39), .A (n_1_40));
OAI22_X1 i_1_122 (.ZN (n_153), .A1 (n_1_811), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_39));
OAI222_X1 i_1_121 (.ZN (n_1_38), .A1 (n_1_874), .A2 (n_1_73), .B1 (n_1_904), .B2 (n_1_72)
    , .C1 (n_1_905), .C2 (n_1_71));
INV_X1 i_1_120 (.ZN (n_1_37), .A (n_1_38));
OAI22_X1 i_1_119 (.ZN (n_152), .A1 (n_1_810), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_37));
OAI222_X1 i_1_118 (.ZN (n_1_36), .A1 (n_1_873), .A2 (n_1_73), .B1 (n_1_903), .B2 (n_1_72)
    , .C1 (n_1_904), .C2 (n_1_71));
INV_X1 i_1_117 (.ZN (n_1_35), .A (n_1_36));
OAI22_X1 i_1_116 (.ZN (n_151), .A1 (n_1_809), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_35));
OAI222_X1 i_1_115 (.ZN (n_1_34), .A1 (n_1_872), .A2 (n_1_73), .B1 (n_1_902), .B2 (n_1_72)
    , .C1 (n_1_903), .C2 (n_1_71));
INV_X1 i_1_114 (.ZN (n_1_33), .A (n_1_34));
OAI22_X1 i_1_113 (.ZN (n_150), .A1 (n_1_808), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_33));
OAI222_X1 i_1_112 (.ZN (n_1_32), .A1 (n_1_871), .A2 (n_1_73), .B1 (n_1_901), .B2 (n_1_72)
    , .C1 (n_1_902), .C2 (n_1_71));
INV_X1 i_1_111 (.ZN (n_1_31), .A (n_1_32));
OAI22_X1 i_1_110 (.ZN (n_149), .A1 (n_1_807), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_31));
OAI222_X1 i_1_109 (.ZN (n_1_30), .A1 (n_1_870), .A2 (n_1_73), .B1 (n_1_900), .B2 (n_1_72)
    , .C1 (n_1_901), .C2 (n_1_71));
INV_X1 i_1_108 (.ZN (n_1_29), .A (n_1_30));
OAI22_X1 i_1_107 (.ZN (n_148), .A1 (n_1_806), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_29));
OAI222_X1 i_1_106 (.ZN (n_1_28), .A1 (n_1_869), .A2 (n_1_73), .B1 (n_1_899), .B2 (n_1_72)
    , .C1 (n_1_900), .C2 (n_1_71));
INV_X1 i_1_105 (.ZN (n_1_27), .A (n_1_28));
OAI22_X1 i_1_104 (.ZN (n_147), .A1 (n_1_805), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_27));
OAI222_X1 i_1_103 (.ZN (n_1_26), .A1 (n_1_868), .A2 (n_1_73), .B1 (n_1_898), .B2 (n_1_72)
    , .C1 (n_1_899), .C2 (n_1_71));
INV_X1 i_1_102 (.ZN (n_1_25), .A (n_1_26));
OAI22_X1 i_1_101 (.ZN (n_146), .A1 (n_1_804), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_25));
OAI222_X1 i_1_100 (.ZN (n_1_24), .A1 (n_1_867), .A2 (n_1_73), .B1 (n_1_897), .B2 (n_1_72)
    , .C1 (n_1_898), .C2 (n_1_71));
INV_X1 i_1_99 (.ZN (n_1_23), .A (n_1_24));
OAI22_X1 i_1_98 (.ZN (n_145), .A1 (n_1_803), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_23));
OAI222_X1 i_1_97 (.ZN (n_1_22), .A1 (n_1_866), .A2 (n_1_73), .B1 (n_1_896), .B2 (n_1_72)
    , .C1 (n_1_897), .C2 (n_1_71));
INV_X1 i_1_96 (.ZN (n_1_21), .A (n_1_22));
OAI22_X1 i_1_95 (.ZN (n_144), .A1 (n_1_802), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_21));
OAI222_X1 i_1_94 (.ZN (n_1_20), .A1 (n_1_865), .A2 (n_1_73), .B1 (n_1_895), .B2 (n_1_72)
    , .C1 (n_1_896), .C2 (n_1_71));
INV_X1 i_1_93 (.ZN (n_1_19), .A (n_1_20));
OAI22_X1 i_1_92 (.ZN (n_143), .A1 (n_1_801), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_19));
OAI222_X1 i_1_91 (.ZN (n_1_18), .A1 (n_1_864), .A2 (n_1_73), .B1 (n_1_894), .B2 (n_1_72)
    , .C1 (n_1_895), .C2 (n_1_71));
INV_X1 i_1_90 (.ZN (n_1_17), .A (n_1_18));
OAI22_X1 i_1_89 (.ZN (n_142), .A1 (n_1_800), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n16), .B2 (n_1_17));
OAI222_X1 i_1_88 (.ZN (n_1_16), .A1 (n_1_863), .A2 (n_1_73), .B1 (n_1_893), .B2 (n_1_72)
    , .C1 (n_1_894), .C2 (n_1_71));
INV_X1 i_1_87 (.ZN (n_1_15), .A (n_1_16));
OAI22_X1 i_1_86 (.ZN (n_141), .A1 (n_1_799), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_15));
OAI222_X1 i_1_85 (.ZN (n_1_14), .A1 (n_1_862), .A2 (n_1_73), .B1 (n_1_892), .B2 (n_1_72)
    , .C1 (n_1_893), .C2 (n_1_71));
INV_X1 i_1_84 (.ZN (n_1_13), .A (n_1_14));
OAI22_X1 i_1_83 (.ZN (n_140), .A1 (n_1_798), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_13));
OAI222_X1 i_1_82 (.ZN (n_1_12), .A1 (n_1_861), .A2 (n_1_73), .B1 (n_1_891), .B2 (n_1_72)
    , .C1 (n_1_892), .C2 (n_1_71));
INV_X1 i_1_81 (.ZN (n_1_11), .A (n_1_12));
OAI22_X1 i_1_80 (.ZN (n_139), .A1 (n_1_797), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_11));
OAI222_X1 i_1_79 (.ZN (n_1_10), .A1 (n_1_860), .A2 (n_1_73), .B1 (n_1_859), .B2 (n_1_72)
    , .C1 (n_1_891), .C2 (n_1_71));
INV_X1 i_1_78 (.ZN (n_1_9), .A (n_1_10));
OAI22_X1 i_1_77 (.ZN (n_138), .A1 (n_1_796), .A2 (hfn_ipo_n13), .B1 (hfn_ipo_n15), .B2 (n_1_9));
NAND3_X1 i_1_76 (.ZN (n_1_8), .A1 (b[0]), .A2 (a[0]), .A3 (hfn_ipo_n13));
OAI21_X1 i_1_75 (.ZN (n_137), .A (n_1_8), .B1 (n_1_795), .B2 (hfn_ipo_n13));
AOI211_X1 i_1_74 (.ZN (n_1_7), .A (reset), .B (resetReg), .C1 (n_1_788), .C2 (n_1_786));
OAI21_X1 i_1_73 (.ZN (n_1_6), .A (n_1_617), .B1 (n_1_922), .B2 (n_1_7));
NOR2_X1 i_1_72 (.ZN (n_136), .A1 (n_1_791), .A2 (n_1_6));
NOR2_X1 i_1_71 (.ZN (n_135), .A1 (n_1_792), .A2 (n_1_6));
NOR2_X1 i_1_70 (.ZN (n_134), .A1 (n_1_793), .A2 (n_1_6));
NOR2_X1 i_1_69 (.ZN (n_133), .A1 (n_1_794), .A2 (n_1_6));
NOR3_X1 i_1_68 (.ZN (n_132), .A1 (\counter[0] ), .A2 (n_267), .A3 (n_1_657));
NOR2_X1 i_1_67 (.ZN (n_131), .A1 (n_1_858), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_66 (.ZN (n_130), .A1 (n_1_857), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_65 (.ZN (n_129), .A1 (n_1_856), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_64 (.ZN (n_128), .A1 (n_1_855), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_63 (.ZN (n_127), .A1 (n_1_854), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_62 (.ZN (n_126), .A1 (n_1_853), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_61 (.ZN (n_125), .A1 (n_1_852), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_60 (.ZN (n_124), .A1 (n_1_851), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_59 (.ZN (n_123), .A1 (n_1_850), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_58 (.ZN (n_122), .A1 (n_1_849), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_57 (.ZN (n_121), .A1 (n_1_848), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_56 (.ZN (n_120), .A1 (n_1_847), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_55 (.ZN (n_119), .A1 (n_1_846), .A2 (n_267));
NOR2_X1 i_1_54 (.ZN (n_118), .A1 (n_1_845), .A2 (n_267));
NOR2_X1 i_1_53 (.ZN (n_117), .A1 (n_1_844), .A2 (n_267));
NOR2_X1 i_1_52 (.ZN (n_116), .A1 (n_1_843), .A2 (n_267));
NOR2_X1 i_1_51 (.ZN (n_115), .A1 (n_1_842), .A2 (n_267));
NOR2_X1 i_1_50 (.ZN (n_114), .A1 (n_1_841), .A2 (n_267));
NOR2_X1 i_1_49 (.ZN (n_113), .A1 (n_1_840), .A2 (n_267));
NOR2_X1 i_1_48 (.ZN (n_112), .A1 (n_1_839), .A2 (n_267));
NOR2_X1 i_1_47 (.ZN (n_111), .A1 (n_1_838), .A2 (n_267));
NOR2_X1 i_1_46 (.ZN (n_110), .A1 (n_1_837), .A2 (n_267));
NOR2_X1 i_1_45 (.ZN (n_109), .A1 (n_1_836), .A2 (n_267));
NOR2_X1 i_1_44 (.ZN (n_108), .A1 (n_1_835), .A2 (n_267));
NOR2_X1 i_1_43 (.ZN (n_107), .A1 (n_1_834), .A2 (n_267));
NOR2_X1 i_1_42 (.ZN (n_106), .A1 (n_1_833), .A2 (n_267));
NOR2_X1 i_1_41 (.ZN (n_105), .A1 (n_1_832), .A2 (n_267));
NOR2_X1 i_1_40 (.ZN (n_104), .A1 (n_1_831), .A2 (n_267));
NOR2_X1 i_1_39 (.ZN (n_103), .A1 (n_1_830), .A2 (n_267));
NOR2_X1 i_1_38 (.ZN (n_102), .A1 (n_1_829), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_37 (.ZN (n_101), .A1 (n_1_828), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_36 (.ZN (n_100), .A1 (n_1_827), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_35 (.ZN (n_99), .A1 (n_1_826), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_34 (.ZN (n_98), .A1 (n_1_825), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_33 (.ZN (n_97), .A1 (n_1_824), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_32 (.ZN (n_96), .A1 (n_1_823), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_31 (.ZN (n_95), .A1 (n_1_822), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_30 (.ZN (n_94), .A1 (n_1_821), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_29 (.ZN (n_93), .A1 (n_1_820), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_28 (.ZN (n_92), .A1 (n_1_819), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_27 (.ZN (n_91), .A1 (n_1_818), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_26 (.ZN (n_90), .A1 (n_1_817), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_25 (.ZN (n_89), .A1 (n_1_816), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_24 (.ZN (n_88), .A1 (n_1_815), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_23 (.ZN (n_87), .A1 (n_1_814), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_22 (.ZN (n_86), .A1 (n_1_813), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_21 (.ZN (n_85), .A1 (n_1_812), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_20 (.ZN (n_84), .A1 (n_1_811), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_19 (.ZN (n_83), .A1 (n_1_810), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_18 (.ZN (n_82), .A1 (n_1_809), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_17 (.ZN (n_81), .A1 (n_1_808), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_16 (.ZN (n_80), .A1 (n_1_807), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_15 (.ZN (n_79), .A1 (n_1_806), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_14 (.ZN (n_78), .A1 (n_1_805), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_13 (.ZN (n_77), .A1 (n_1_804), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_12 (.ZN (n_76), .A1 (n_1_803), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_11 (.ZN (n_75), .A1 (n_1_802), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_10 (.ZN (n_74), .A1 (n_1_801), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_9 (.ZN (n_73), .A1 (n_1_800), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_8 (.ZN (n_72), .A1 (n_1_799), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_7 (.ZN (n_71), .A1 (n_1_798), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_6 (.ZN (n_70), .A1 (n_1_797), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_5 (.ZN (n_69), .A1 (n_1_796), .A2 (hfn_ipo_n17));
NOR2_X1 i_1_4 (.ZN (n_68), .A1 (n_1_795), .A2 (hfn_ipo_n17));
AND2_X1 i_1_3 (.ZN (n_67), .A1 (en), .A2 (reset));
HA_X1 i_1_2 (.CO (n_1_2), .S (n_1_5), .A (\counter[3] ), .B (n_1_1));
HA_X1 i_1_1 (.CO (n_1_1), .S (n_1_4), .A (\counter[2] ), .B (n_1_0));
HA_X1 i_1_0 (.CO (n_1_0), .S (n_1_3), .A (\counter[1] ), .B (\counter[0] ));
datapath__0_74 i_41 (.p_1 ({n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, 
    n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, 
    n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, 
    n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, 
    n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
    n_4, n_3}), .aux ({\aux[63] , \aux[62] , \aux[61] , \aux[60] , \aux[59] , \aux[58] , 
    \aux[57] , \aux[56] , \aux[55] , \aux[54] , \aux[53] , \aux[52] , \aux[51] , 
    \aux[50] , \aux[49] , \aux[48] , \aux[47] , \aux[46] , \aux[45] , \aux[44] , 
    \aux[43] , \aux[42] , \aux[41] , \aux[40] , \aux[39] , \aux[38] , \aux[37] , 
    \aux[36] , \aux[35] , \aux[34] , \aux[33] , \aux[32] , \aux[31] , \aux[30] , 
    \aux[29] , \aux[28] , \aux[27] , \aux[26] , \aux[25] , \aux[24] , \aux[23] , 
    \aux[22] , \aux[21] , \aux[20] , \aux[19] , \aux[18] , \aux[17] , \aux[16] , 
    \aux[15] , \aux[14] , \aux[13] , \aux[12] , \aux[11] , \aux[10] , \aux[9] , \aux[8] , 
    \aux[7] , \aux[6] , \aux[5] , \aux[4] , \aux[3] , \aux[2] , \aux[1] , \aux[0] })
    , .p_0 ({n_264, n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, 
    n_254, n_253, n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, 
    n_243, n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, 
    n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, n_222, 
    n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, 
    n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201}));
DFF_X1 enableOutput_reg (.Q (enableOutput), .CK (CTS_n_tid0_153), .D (n_268));
datapath i_0 (.firstInputComplement ({\firstInputComplement[31] , \firstInputComplement[30] , 
    \firstInputComplement[29] , \firstInputComplement[28] , \firstInputComplement[27] , 
    \firstInputComplement[26] , \firstInputComplement[25] , \firstInputComplement[24] , 
    \firstInputComplement[23] , \firstInputComplement[22] , \firstInputComplement[21] , 
    \firstInputComplement[20] , \firstInputComplement[19] , \firstInputComplement[18] , 
    \firstInputComplement[17] , \firstInputComplement[16] , \firstInputComplement[15] , 
    \firstInputComplement[14] , \firstInputComplement[13] , \firstInputComplement[12] , 
    \firstInputComplement[11] , \firstInputComplement[10] , \firstInputComplement[9] , 
    \firstInputComplement[8] , \firstInputComplement[7] , \firstInputComplement[6] , 
    \firstInputComplement[5] , \firstInputComplement[4] , \firstInputComplement[3] , 
    \firstInputComplement[2] , \firstInputComplement[1] , uc_0}), .a ({a[31], a[30], 
    a[29], a[28], a[27], a[26], a[25], a[24], a[23], a[22], a[21], a[20], a[19], 
    a[18], a[17], a[16], a[15], a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7], 
    a[6], a[5], a[4], a[3], a[2], a[1], a[0]}));
BUF_X8 hfn_ipo_c17 (.Z (hfn_ipo_n17), .A (n_267));
INV_X16 CTS_L6_c_tid0_72 (.ZN (CTS_n_tid0_82), .A (CTS_n_tid0_84));
BUF_X2 hfn_ipo_c15 (.Z (hfn_ipo_n15), .A (n_1_785));
BUF_X2 hfn_ipo_c16 (.Z (hfn_ipo_n16), .A (n_1_785));
BUF_X8 hfn_ipo_c13 (.Z (hfn_ipo_n13), .A (n_1_784));
BUF_X8 hfn_ipo_c14 (.Z (hfn_ipo_n14), .A (n_1_784));
BUF_X1 drc_ipo_c19 (.Z (drc_ipo_n19), .A (n_1_665));
INV_X8 CTS_L7_c_tid0_71 (.ZN (CTS_n_tid0_81), .A (CTS_n_tid0_82));
INV_X4 CTS_L5_c_tid0_154 (.ZN (clk_CTS_0_PP_8), .A (CTS_n_tid0_247));
INV_X4 CTS_L6_c_tid0_126 (.ZN (CTS_n_tid0_153), .A (clk_CTS_0_PP_8));
BUF_X16 CTS_L8_c_tid1_67 (.Z (CTS_n_tid1_76), .A (CTS_n_tid1_73));
INV_X4 CTS_L6_c_tid0_141 (.ZN (CTS_n_tid0_189), .A (CTS_n_tid0_206));
INV_X16 CTS_L5_c_tid0_153 (.ZN (CTS_n_tid0_206), .A (CTS_n_tid0_247));
BUF_X1 CLOCK_sgo__c183 (.Z (CLOCK_sgo__n273), .A (n_1_640));
BUF_X8 CTS_L4_c_tid0_181 (.Z (CTS_n_tid0_247), .A (clk_CTS_0_PP_14));

endmodule //radix4Booth

module registerNbits__0_87 (clk_CTS_0_PP_0, clk_CTS_0_PP_1, clk, reset, en, inp, 
    out);

output [31:0] out;
output clk_CTS_0_PP_0;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_1;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid0_6;
wire CLOCK_slh__n49;
wire CLOCK_slh__n51;
wire CLOCK_slh__n53;
wire CLOCK_slh__n55;
wire CLOCK_slh__n57;
wire CLOCK_slh__n59;
wire CLOCK_slh__n61;
wire CLOCK_slh__n63;
wire CLOCK_slh__n65;
wire CLOCK_slh__n67;
wire CLOCK_slh__n69;
wire CLOCK_slh__n71;
wire CLOCK_slh__n73;
wire CLOCK_slh__n75;
wire CLOCK_slh__n77;
wire CLOCK_slh__n79;
wire CLOCK_slh__n81;
wire CLOCK_slh__n83;
wire CLOCK_slh__n85;
wire CLOCK_slh__n87;
wire CLOCK_slh__n89;
wire CLOCK_slh__n90;
wire CLOCK_slh__n91;
wire CLOCK_slh__n92;
wire CLOCK_slh__n93;
wire CLOCK_slh__n94;
wire CLOCK_slh__n95;
wire CLOCK_slh__n96;
wire CLOCK_slh__n97;
wire CLOCK_slh__n98;
wire CLOCK_slh__n99;
wire CLOCK_slh__n100;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n95), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n91), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n71), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n83), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n97), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n90), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n63), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n81), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n100), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n61), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n79), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n67), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n94), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n49), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n59), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n57), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n96), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n85), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n77), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n73), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n93), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n92), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n69), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n89), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n87), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n65), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n99), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n75), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n98), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n53), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n51), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n55), .A1 (n_0_0), .A2 (inp[0]));
INV_X2 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
INV_X4 CTS_L3_c_tid0_7 (.ZN (clk_CTS_0_PP_0), .A (CTS_n_tid0_6));
INV_X4 CTS_L2_c_tid0_8 (.ZN (CTS_n_tid0_6), .A (clk_CTS_0_PP_1));
CLKBUF_X1 CLOCK_slh__c22 (.Z (n_20), .A (CLOCK_slh__n49));
CLKBUF_X1 CLOCK_slh__c24 (.Z (n_3), .A (CLOCK_slh__n51));
CLKBUF_X1 CLOCK_slh__c26 (.Z (n_4), .A (CLOCK_slh__n53));
CLKBUF_X1 CLOCK_slh__c28 (.Z (n_2), .A (CLOCK_slh__n55));
CLKBUF_X1 CLOCK_slh__c30 (.Z (n_18), .A (CLOCK_slh__n57));
CLKBUF_X1 CLOCK_slh__c32 (.Z (n_19), .A (CLOCK_slh__n59));
CLKBUF_X1 CLOCK_slh__c34 (.Z (n_24), .A (CLOCK_slh__n61));
CLKBUF_X1 CLOCK_slh__c36 (.Z (n_27), .A (CLOCK_slh__n63));
CLKBUF_X1 CLOCK_slh__c38 (.Z (n_8), .A (CLOCK_slh__n65));
CLKBUF_X1 CLOCK_slh__c40 (.Z (n_22), .A (CLOCK_slh__n67));
CLKBUF_X1 CLOCK_slh__c42 (.Z (n_11), .A (CLOCK_slh__n69));
CLKBUF_X1 CLOCK_slh__c44 (.Z (n_31), .A (CLOCK_slh__n71));
CLKBUF_X1 CLOCK_slh__c46 (.Z (n_14), .A (CLOCK_slh__n73));
CLKBUF_X1 CLOCK_slh__c48 (.Z (n_6), .A (CLOCK_slh__n75));
CLKBUF_X1 CLOCK_slh__c50 (.Z (n_15), .A (CLOCK_slh__n77));
CLKBUF_X1 CLOCK_slh__c52 (.Z (n_23), .A (CLOCK_slh__n79));
CLKBUF_X1 CLOCK_slh__c54 (.Z (n_26), .A (CLOCK_slh__n81));
CLKBUF_X1 CLOCK_slh__c56 (.Z (n_30), .A (CLOCK_slh__n83));
CLKBUF_X1 CLOCK_slh__c58 (.Z (n_16), .A (CLOCK_slh__n85));
CLKBUF_X1 CLOCK_slh__c60 (.Z (n_9), .A (CLOCK_slh__n87));
CLKBUF_X1 CLOCK_slh__c62 (.Z (n_10), .A (CLOCK_slh__n89));
CLKBUF_X1 CLOCK_slh__c63 (.Z (n_28), .A (CLOCK_slh__n90));
CLKBUF_X1 CLOCK_slh__c64 (.Z (n_32), .A (CLOCK_slh__n91));
CLKBUF_X1 CLOCK_slh__c65 (.Z (n_12), .A (CLOCK_slh__n92));
CLKBUF_X1 CLOCK_slh__c66 (.Z (n_13), .A (CLOCK_slh__n93));
CLKBUF_X1 CLOCK_slh__c67 (.Z (n_21), .A (CLOCK_slh__n94));
CLKBUF_X1 CLOCK_slh__c68 (.Z (n_33), .A (CLOCK_slh__n95));
CLKBUF_X1 CLOCK_slh__c69 (.Z (n_17), .A (CLOCK_slh__n96));
CLKBUF_X1 CLOCK_slh__c70 (.Z (n_29), .A (CLOCK_slh__n97));
CLKBUF_X1 CLOCK_slh__c71 (.Z (n_5), .A (CLOCK_slh__n98));
CLKBUF_X1 CLOCK_slh__c72 (.Z (n_7), .A (CLOCK_slh__n99));
CLKBUF_X1 CLOCK_slh__c73 (.Z (n_25), .A (CLOCK_slh__n100));

endmodule //registerNbits__0_87

module registerNbits__0_84 (clk_CTS_0_PP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CLOCK_slh__n20;
wire CLOCK_slh__n22;
wire CLOCK_slh__n24;
wire CLOCK_slh__n26;
wire CLOCK_slh__n28;
wire CLOCK_slh__n30;
wire CLOCK_slh__n32;
wire CLOCK_slh__n34;
wire CLOCK_slh__n36;
wire CLOCK_slh__n38;
wire CLOCK_slh__n40;
wire CLOCK_slh__n42;
wire CLOCK_slh__n44;
wire CLOCK_slh__n46;
wire CLOCK_slh__n48;
wire CLOCK_slh__n50;
wire CLOCK_slh__n52;
wire CLOCK_slh__n54;
wire CLOCK_slh__n56;
wire CLOCK_slh__n58;
wire CLOCK_slh__n60;
wire CLOCK_slh__n62;
wire CLOCK_slh__n64;
wire CLOCK_slh__n66;
wire CLOCK_slh__n68;
wire CLOCK_slh__n70;
wire CLOCK_slh__n72;
wire CLOCK_slh__n74;
wire CLOCK_slh__n76;
wire CLOCK_slh__n78;
wire CLOCK_slh__n80;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n44), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n42), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n60), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n40), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n72), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n78), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n46), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n76), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n56), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n74), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n80), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n66), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n70), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n64), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n68), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n58), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n62), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n34), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n50), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n24), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n32), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n48), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n54), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n22), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n30), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n20), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n26), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n28), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n36), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n38), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n52), .A1 (n_0_0), .A2 (inp[0]));
INV_X2 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X1 CLOCK_slh__c7 (.Z (n_7), .A (CLOCK_slh__n20));
CLKBUF_X1 CLOCK_slh__c9 (.Z (n_9), .A (CLOCK_slh__n22));
CLKBUF_X1 CLOCK_slh__c11 (.Z (n_13), .A (CLOCK_slh__n24));
CLKBUF_X1 CLOCK_slh__c13 (.Z (n_6), .A (CLOCK_slh__n26));
CLKBUF_X1 CLOCK_slh__c15 (.Z (n_5), .A (CLOCK_slh__n28));
CLKBUF_X1 CLOCK_slh__c17 (.Z (n_8), .A (CLOCK_slh__n30));
CLKBUF_X1 CLOCK_slh__c19 (.Z (n_12), .A (CLOCK_slh__n32));
CLKBUF_X1 CLOCK_slh__c21 (.Z (n_15), .A (CLOCK_slh__n34));
CLKBUF_X1 CLOCK_slh__c23 (.Z (n_4), .A (CLOCK_slh__n36));
CLKBUF_X1 CLOCK_slh__c25 (.Z (n_3), .A (CLOCK_slh__n38));
CLKBUF_X1 CLOCK_slh__c27 (.Z (n_30), .A (CLOCK_slh__n40));
CLKBUF_X1 CLOCK_slh__c29 (.Z (n_32), .A (CLOCK_slh__n42));
CLKBUF_X1 CLOCK_slh__c31 (.Z (n_33), .A (CLOCK_slh__n44));
CLKBUF_X1 CLOCK_slh__c33 (.Z (n_27), .A (CLOCK_slh__n46));
CLKBUF_X1 CLOCK_slh__c35 (.Z (n_11), .A (CLOCK_slh__n48));
CLKBUF_X1 CLOCK_slh__c37 (.Z (n_14), .A (CLOCK_slh__n50));
CLKBUF_X1 CLOCK_slh__c39 (.Z (n_2), .A (CLOCK_slh__n52));
CLKBUF_X1 CLOCK_slh__c41 (.Z (n_10), .A (CLOCK_slh__n54));
CLKBUF_X1 CLOCK_slh__c43 (.Z (n_25), .A (CLOCK_slh__n56));
CLKBUF_X1 CLOCK_slh__c45 (.Z (n_17), .A (CLOCK_slh__n58));
CLKBUF_X1 CLOCK_slh__c47 (.Z (n_31), .A (CLOCK_slh__n60));
CLKBUF_X1 CLOCK_slh__c49 (.Z (n_16), .A (CLOCK_slh__n62));
CLKBUF_X1 CLOCK_slh__c51 (.Z (n_19), .A (CLOCK_slh__n64));
CLKBUF_X1 CLOCK_slh__c53 (.Z (n_22), .A (CLOCK_slh__n66));
CLKBUF_X1 CLOCK_slh__c55 (.Z (n_18), .A (CLOCK_slh__n68));
CLKBUF_X1 CLOCK_slh__c57 (.Z (n_21), .A (CLOCK_slh__n70));
CLKBUF_X1 CLOCK_slh__c59 (.Z (n_29), .A (CLOCK_slh__n72));
CLKBUF_X1 CLOCK_slh__c61 (.Z (n_24), .A (CLOCK_slh__n74));
CLKBUF_X1 CLOCK_slh__c63 (.Z (n_26), .A (CLOCK_slh__n76));
CLKBUF_X1 CLOCK_slh__c65 (.Z (n_28), .A (CLOCK_slh__n78));
CLKBUF_X1 CLOCK_slh__c67 (.Z (n_23), .A (CLOCK_slh__n80));

endmodule //registerNbits__0_84

module integrationMult (inputA, inputB, clk, reset, en, result);

output [63:0] result;
input clk;
input en;
input [31:0] inputA;
input [31:0] inputB;
input reset;
wire CTS_n_tid0_24;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire enableOutput;
wire \outB_reg[31] ;
wire \outB_reg[30] ;
wire \outB_reg[29] ;
wire \outB_reg[28] ;
wire \outB_reg[27] ;
wire \outB_reg[26] ;
wire \outB_reg[25] ;
wire \outB_reg[24] ;
wire \outB_reg[23] ;
wire \outB_reg[22] ;
wire \outB_reg[21] ;
wire \outB_reg[20] ;
wire \outB_reg[19] ;
wire \outB_reg[18] ;
wire \outB_reg[17] ;
wire \outB_reg[16] ;
wire \outB_reg[15] ;
wire \outB_reg[14] ;
wire \outB_reg[13] ;
wire \outB_reg[12] ;
wire \outB_reg[11] ;
wire \outB_reg[10] ;
wire \outB_reg[9] ;
wire \outB_reg[8] ;
wire \outB_reg[7] ;
wire \outB_reg[6] ;
wire \outB_reg[5] ;
wire \outB_reg[4] ;
wire \outB_reg[3] ;
wire \outB_reg[2] ;
wire \outB_reg[1] ;
wire \outB_reg[0] ;
wire \outA_reg[31] ;
wire \outA_reg[30] ;
wire \outA_reg[29] ;
wire \outA_reg[28] ;
wire \outA_reg[27] ;
wire \outA_reg[26] ;
wire \outA_reg[25] ;
wire \outA_reg[24] ;
wire \outA_reg[23] ;
wire \outA_reg[22] ;
wire \outA_reg[21] ;
wire \outA_reg[20] ;
wire \outA_reg[19] ;
wire \outA_reg[18] ;
wire \outA_reg[17] ;
wire \outA_reg[16] ;
wire \outA_reg[15] ;
wire \outA_reg[14] ;
wire \outA_reg[13] ;
wire \outA_reg[12] ;
wire \outA_reg[11] ;
wire \outA_reg[10] ;
wire \outA_reg[9] ;
wire \outA_reg[8] ;
wire \outA_reg[7] ;
wire \outA_reg[6] ;
wire \outA_reg[5] ;
wire \outA_reg[4] ;
wire \outA_reg[3] ;
wire \outA_reg[2] ;
wire \outA_reg[1] ;
wire \outA_reg[0] ;
wire CLOCK_n_tid0_127;
wire CTS_n_tid0_42;


registerNbits outA (.out ({result[31], result[30], result[29], result[28], result[27], 
    result[26], result[25], result[24], result[23], result[22], result[21], result[20], 
    result[19], result[18], result[17], result[16], result[15], result[14], result[13], 
    result[12], result[11], result[10], result[9], result[8], result[7], result[6], 
    result[5], result[4], result[3], result[2], result[1], result[0]}), .en (enableOutput)
    , .inp ({\outB_reg[31] , \outB_reg[30] , \outB_reg[29] , \outB_reg[28] , \outB_reg[27] , 
    \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , \outB_reg[23] , \outB_reg[22] , 
    \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , \outB_reg[18] , \outB_reg[17] , 
    \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , \outB_reg[13] , \outB_reg[12] , 
    \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , \outB_reg[8] , \outB_reg[7] , 
    \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , 
    \outB_reg[0] }), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_42));
registerNbits__0_90 outB (.out ({result[63], result[62], result[61], result[60], 
    result[59], result[58], result[57], result[56], result[55], result[54], result[53], 
    result[52], result[51], result[50], result[49], result[48], result[47], result[46], 
    result[45], result[44], result[43], result[42], result[41], result[40], result[39], 
    result[38], result[37], result[36], result[35], result[34], result[33], result[32]})
    , .en (enableOutput), .inp ({\outA_reg[31] , \outA_reg[30] , \outA_reg[29] , 
    \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , \outA_reg[24] , 
    \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , \outA_reg[19] , 
    \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , \outA_reg[14] , 
    \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , \outA_reg[9] , 
    \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , 
    \outA_reg[2] , \outA_reg[1] , \outA_reg[0] }), .reset (reset), .clk_CTS_0_PP_8 (CTS_n_tid0_24));
radix4Booth radix4BoothIns (.enableOutput (enableOutput), .result ({\outA_reg[31] , 
    \outA_reg[30] , \outA_reg[29] , \outA_reg[28] , \outA_reg[27] , \outA_reg[26] , 
    \outA_reg[25] , \outA_reg[24] , \outA_reg[23] , \outA_reg[22] , \outA_reg[21] , 
    \outA_reg[20] , \outA_reg[19] , \outA_reg[18] , \outA_reg[17] , \outA_reg[16] , 
    \outA_reg[15] , \outA_reg[14] , \outA_reg[13] , \outA_reg[12] , \outA_reg[11] , 
    \outA_reg[10] , \outA_reg[9] , \outA_reg[8] , \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , 
    \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , \outA_reg[1] , \outA_reg[0] , \outB_reg[31] , 
    \outB_reg[30] , \outB_reg[29] , \outB_reg[28] , \outB_reg[27] , \outB_reg[26] , 
    \outB_reg[25] , \outB_reg[24] , \outB_reg[23] , \outB_reg[22] , \outB_reg[21] , 
    \outB_reg[20] , \outB_reg[19] , \outB_reg[18] , \outB_reg[17] , \outB_reg[16] , 
    \outB_reg[15] , \outB_reg[14] , \outB_reg[13] , \outB_reg[12] , \outB_reg[11] , 
    \outB_reg[10] , \outB_reg[9] , \outB_reg[8] , \outB_reg[7] , \outB_reg[6] , \outB_reg[5] , 
    \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , \outB_reg[0] }), .clk_CTS_0_PP_8 (CTS_n_tid0_24)
    , .a ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , \A_reg[27] , \A_reg[26] , 
    \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , \A_reg[21] , \A_reg[20] , 
    \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , \A_reg[15] , \A_reg[14] , 
    \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , \A_reg[9] , \A_reg[8] , \A_reg[7] , 
    \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , \A_reg[1] , \A_reg[0] })
    , .b ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , \B_reg[26] , 
    \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , \B_reg[20] , 
    \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , \B_reg[14] , 
    \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , \B_reg[8] , \B_reg[7] , 
    \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] })
    , .en (en), .reset (reset), .clk_CTS_0_PP_14 (CTS_n_tid0_42));
registerNbits__0_87 regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , 
    \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , 
    \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , 
    \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , 
    \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .clk_CTS_0_PP_0 (CTS_n_tid0_42), .en (en)
    , .inp ({inputB[31], inputB[30], inputB[29], inputB[28], inputB[27], inputB[26], 
    inputB[25], inputB[24], inputB[23], inputB[22], inputB[21], inputB[20], inputB[19], 
    inputB[18], inputB[17], inputB[16], inputB[15], inputB[14], inputB[13], inputB[12], 
    inputB[11], inputB[10], inputB[9], inputB[8], inputB[7], inputB[6], inputB[5], 
    inputB[4], inputB[3], inputB[2], inputB[1], inputB[0]}), .reset (reset), .clk_CTS_0_PP_1 (CLOCK_n_tid0_127));
registerNbits__0_84 regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .en (en), .inp ({inputA[31], inputA[30], 
    inputA[29], inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], 
    inputA[22], inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], 
    inputA[15], inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], 
    inputA[8], inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], 
    inputA[1], inputA[0]}), .reset (reset), .clk_CTS_0_PP_0 (CTS_n_tid0_42));
BUF_X8 CTS_L1_tid0__c1_tid0__c63 (.Z (CLOCK_n_tid0_127), .A (clk));

endmodule //integrationMult


